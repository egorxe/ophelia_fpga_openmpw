VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_ctrl
  CLASS BLOCK ;
  FOREIGN efuse_ctrl ;
  ORIGIN 0.000 0.000 ;
  SIZE 2175.000 BY 2350.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 25.920 15.380 27.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 15.380 217.520 29.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 768.115 217.520 789.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 1528.115 217.520 1549.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 2288.115 217.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 15.380 407.520 32.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 767.505 407.520 792.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 1527.505 407.520 1552.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 2287.505 407.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 15.380 597.520 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 767.505 597.520 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 1527.505 597.520 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 2287.505 597.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 15.380 787.520 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 767.530 787.520 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 1527.530 787.520 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 2287.530 787.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 15.380 977.520 32.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 767.505 977.520 792.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 1527.505 977.520 1552.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 2287.505 977.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1165.920 15.380 1167.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1355.920 15.380 1357.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 15.380 1547.520 29.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 767.530 1547.520 789.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 1527.530 1547.520 1549.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 2287.530 1547.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 15.380 1737.520 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 767.505 1737.520 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 1527.505 1737.520 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 2287.505 1737.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 15.380 1927.520 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 767.505 1927.520 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 1527.505 1927.520 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 2287.505 1927.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 15.380 2117.520 32.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 767.530 2117.520 792.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 1527.530 2117.520 1552.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 2287.530 2117.520 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 23.220 111.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 783.700 199.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 1544.180 287.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 783.700 111.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 23.220 199.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 1544.180 375.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 1544.180 111.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 23.220 287.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 783.700 375.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 1544.180 199.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 783.700 287.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 23.220 375.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.040 23.220 463.640 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.960 783.700 551.560 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 1544.180 640.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.040 783.700 463.640 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.960 23.220 551.560 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 1544.180 727.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.040 1544.180 463.640 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 23.220 640.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 783.700 727.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.960 1544.180 551.560 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 783.700 640.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 23.220 727.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 23.220 815.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 783.700 903.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 990.120 1544.180 991.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 783.700 815.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 23.220 903.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.040 1544.180 1079.640 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 1544.180 815.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 990.120 23.220 991.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.040 783.700 1079.640 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 1544.180 903.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 990.120 783.700 991.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.040 23.220 1079.640 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 23.220 1256.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 1544.180 1431.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 783.700 1256.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 1544.180 1519.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 1544.180 1256.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 23.220 1431.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 783.700 1519.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 783.700 1431.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 23.220 1519.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 23.220 1607.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.040 783.700 1695.640 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1781.960 1544.180 1783.560 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 783.700 1607.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.040 23.220 1695.640 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 1544.180 1872.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 1544.180 1607.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1781.960 23.220 1783.560 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 783.700 1872.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.040 1544.180 1695.640 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1781.960 783.700 1783.560 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 23.220 1872.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 23.220 1959.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 783.700 2047.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2143.720 1544.180 2145.320 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 783.700 1959.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 23.220 2047.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 1544.180 1959.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2143.720 23.220 2145.320 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 1544.180 2047.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2143.720 783.700 2145.320 1533.020 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 35.520 15.380 37.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 15.380 227.120 29.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 767.530 227.120 789.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 1527.530 227.120 1549.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 2287.530 227.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 15.380 417.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 767.505 417.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 1527.505 417.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 2287.505 417.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 15.380 607.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 767.505 607.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 1527.505 607.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 2287.505 607.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 15.380 797.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 767.530 797.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 1527.530 797.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 2287.530 797.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 985.520 15.380 987.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1175.520 15.380 1177.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 15.380 1367.120 29.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 767.530 1367.120 789.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 1527.530 1367.120 1549.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 2287.530 1367.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 15.380 1557.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 767.505 1557.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 1527.505 1557.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 2287.505 1557.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 15.380 1747.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 767.505 1747.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 1527.505 1747.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 2287.505 1747.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 15.380 1937.120 32.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 767.530 1937.120 792.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 1527.530 1937.120 1552.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 2287.530 1937.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 15.380 2127.120 30.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 768.115 2127.120 790.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 1528.115 2127.120 1550.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 2288.115 2127.120 2332.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 23.220 122.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 783.700 209.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 1544.180 297.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 783.700 122.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 23.220 209.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 1544.180 385.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 1544.180 122.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 23.220 297.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 783.700 385.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 1544.180 209.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 783.700 297.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 23.220 385.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.120 23.220 473.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.040 783.700 561.640 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 1544.180 650.120 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.120 783.700 473.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.040 23.220 561.640 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 1544.180 738.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.120 1544.180 473.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 23.220 650.120 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 783.700 738.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.040 1544.180 561.640 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 783.700 650.120 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 23.220 738.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 23.220 825.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 783.700 913.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1000.200 1544.180 1001.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 783.700 825.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 23.220 913.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.120 1544.180 1089.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 1544.180 825.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1000.200 23.220 1001.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.120 783.700 1089.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 1544.180 913.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1000.200 783.700 1001.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.120 23.220 1089.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 23.220 1266.120 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1347.400 783.700 1349.000 1529.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 1544.180 1441.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 783.700 1266.120 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1347.400 23.220 1349.000 768.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 1544.180 1529.880 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 1544.180 1266.120 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 23.220 1441.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 783.700 1529.880 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1347.400 1544.180 1349.000 2289.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 783.700 1441.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 23.220 1529.880 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 23.220 1617.800 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.120 783.700 1705.720 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.040 1544.180 1793.640 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 783.700 1617.800 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.120 23.220 1705.720 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 1544.180 1882.120 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 1544.180 1617.800 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.040 23.220 1793.640 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 783.700 1882.120 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.120 1544.180 1705.720 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.040 783.700 1793.640 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 23.220 1882.120 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 23.220 1970.040 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 783.700 2057.960 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2153.800 1544.180 2155.400 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 783.700 1970.040 1533.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 23.220 2057.960 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 1544.180 1970.040 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2153.800 23.220 2155.400 772.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 1544.180 2057.960 2293.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2153.800 783.700 2155.400 1533.020 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 547.680 4.000 548.240 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 2346.000 2040.080 2349.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1.000 1095.920 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 2346.000 665.840 2349.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 823.200 4.000 823.760 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 840.000 2174.000 840.560 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1216.320 2346.000 1216.880 2349.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 16.800 2174.000 17.360 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 1391.040 2174.000 1391.600 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1918.560 1.000 1919.120 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 1663.200 2174.000 1663.760 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 272.160 4.000 272.720 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1488.480 2346.000 1489.040 2349.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 2346.000 1764.560 2349.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1646.400 4.000 1646.960 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 2346.000 390.320 2349.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1646.400 1.000 1646.960 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1918.560 4.000 1919.120 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 292.320 2174.000 292.880 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 1.000 272.720 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 1.000 548.240 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 2346.000 118.160 2349.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 564.480 2174.000 565.040 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 1.000 823.760 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 1938.720 2174.000 1939.280 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 2214.240 2174.000 2214.800 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1370.880 4.000 1371.440 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 2346.000 941.360 2349.000 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1370.880 1.000 1371.440 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1095.360 4.000 1095.920 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2194.080 4.000 2194.640 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2171.000 1115.520 2174.000 1116.080 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2167.760 2332.700 ;
      LAYER Metal2 ;
        RECT 8.540 2345.700 117.300 2346.000 ;
        RECT 118.460 2345.700 389.460 2346.000 ;
        RECT 390.620 2345.700 664.980 2346.000 ;
        RECT 666.140 2345.700 940.500 2346.000 ;
        RECT 941.660 2345.700 1216.020 2346.000 ;
        RECT 1217.180 2345.700 1488.180 2346.000 ;
        RECT 1489.340 2345.700 1763.700 2346.000 ;
        RECT 1764.860 2345.700 2039.220 2346.000 ;
        RECT 2040.380 2345.700 2165.380 2346.000 ;
        RECT 8.540 4.300 2165.380 2345.700 ;
        RECT 8.540 1.770 271.860 4.300 ;
        RECT 273.020 1.770 547.380 4.300 ;
        RECT 548.540 1.770 822.900 4.300 ;
        RECT 824.060 1.770 1095.060 4.300 ;
        RECT 1096.220 1.770 1370.580 4.300 ;
        RECT 1371.740 1.770 1646.100 4.300 ;
        RECT 1647.260 1.770 1918.260 4.300 ;
        RECT 1919.420 1.770 2165.380 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 2215.100 2171.000 2332.540 ;
        RECT 4.000 2213.940 2170.700 2215.100 ;
        RECT 4.000 2194.940 2171.000 2213.940 ;
        RECT 4.300 2193.780 2171.000 2194.940 ;
        RECT 4.000 1939.580 2171.000 2193.780 ;
        RECT 4.000 1938.420 2170.700 1939.580 ;
        RECT 4.000 1919.420 2171.000 1938.420 ;
        RECT 4.300 1918.260 2171.000 1919.420 ;
        RECT 4.000 1664.060 2171.000 1918.260 ;
        RECT 4.000 1662.900 2170.700 1664.060 ;
        RECT 4.000 1647.260 2171.000 1662.900 ;
        RECT 4.300 1646.100 2171.000 1647.260 ;
        RECT 4.000 1391.900 2171.000 1646.100 ;
        RECT 4.000 1390.740 2170.700 1391.900 ;
        RECT 4.000 1371.740 2171.000 1390.740 ;
        RECT 4.300 1370.580 2171.000 1371.740 ;
        RECT 4.000 1116.380 2171.000 1370.580 ;
        RECT 4.000 1115.220 2170.700 1116.380 ;
        RECT 4.000 1096.220 2171.000 1115.220 ;
        RECT 4.300 1095.060 2171.000 1096.220 ;
        RECT 4.000 840.860 2171.000 1095.060 ;
        RECT 4.000 839.700 2170.700 840.860 ;
        RECT 4.000 824.060 2171.000 839.700 ;
        RECT 4.300 822.900 2171.000 824.060 ;
        RECT 4.000 565.340 2171.000 822.900 ;
        RECT 4.000 564.180 2170.700 565.340 ;
        RECT 4.000 548.540 2171.000 564.180 ;
        RECT 4.300 547.380 2171.000 548.540 ;
        RECT 4.000 293.180 2171.000 547.380 ;
        RECT 4.000 292.020 2170.700 293.180 ;
        RECT 4.000 273.020 2171.000 292.020 ;
        RECT 4.300 271.860 2171.000 273.020 ;
        RECT 4.000 17.660 2171.000 271.860 ;
        RECT 4.000 16.500 2170.700 17.660 ;
        RECT 4.000 1.260 2171.000 16.500 ;
      LAYER Metal4 ;
        RECT 16.940 15.080 25.620 2330.070 ;
        RECT 27.820 15.080 35.220 2330.070 ;
        RECT 37.420 2293.800 215.620 2330.070 ;
        RECT 37.420 1543.880 110.060 2293.800 ;
        RECT 112.260 1543.880 120.140 2293.800 ;
        RECT 122.340 1543.880 197.980 2293.800 ;
        RECT 200.180 1543.880 208.060 2293.800 ;
        RECT 210.260 2287.815 215.620 2293.800 ;
        RECT 217.820 2287.815 225.220 2330.070 ;
        RECT 210.260 2287.230 225.220 2287.815 ;
        RECT 227.420 2293.800 405.620 2330.070 ;
        RECT 227.420 2287.230 285.900 2293.800 ;
        RECT 210.260 1550.020 285.900 2287.230 ;
        RECT 210.260 1543.880 215.620 1550.020 ;
        RECT 37.420 1533.320 215.620 1543.880 ;
        RECT 37.420 783.400 110.060 1533.320 ;
        RECT 112.260 783.400 120.140 1533.320 ;
        RECT 122.340 783.400 197.980 1533.320 ;
        RECT 200.180 783.400 208.060 1533.320 ;
        RECT 210.260 1527.815 215.620 1533.320 ;
        RECT 217.820 1527.815 225.220 1550.020 ;
        RECT 210.260 1527.230 225.220 1527.815 ;
        RECT 227.420 1543.880 285.900 1550.020 ;
        RECT 288.100 1543.880 295.980 2293.800 ;
        RECT 298.180 1543.880 373.820 2293.800 ;
        RECT 376.020 1543.880 383.900 2293.800 ;
        RECT 386.100 2287.205 405.620 2293.800 ;
        RECT 407.820 2287.205 415.220 2330.070 ;
        RECT 417.420 2293.800 595.620 2330.070 ;
        RECT 417.420 2287.205 461.740 2293.800 ;
        RECT 386.100 1552.570 461.740 2287.205 ;
        RECT 386.100 1552.545 415.220 1552.570 ;
        RECT 386.100 1543.880 405.620 1552.545 ;
        RECT 227.420 1533.320 405.620 1543.880 ;
        RECT 227.420 1527.230 285.900 1533.320 ;
        RECT 210.260 790.020 285.900 1527.230 ;
        RECT 210.260 783.400 215.620 790.020 ;
        RECT 37.420 772.840 215.620 783.400 ;
        RECT 37.420 22.920 110.060 772.840 ;
        RECT 112.260 22.920 120.140 772.840 ;
        RECT 122.340 22.920 197.980 772.840 ;
        RECT 200.180 22.920 208.060 772.840 ;
        RECT 210.260 767.815 215.620 772.840 ;
        RECT 217.820 767.815 225.220 790.020 ;
        RECT 210.260 767.230 225.220 767.815 ;
        RECT 227.420 783.400 285.900 790.020 ;
        RECT 288.100 783.400 295.980 1533.320 ;
        RECT 298.180 783.400 373.820 1533.320 ;
        RECT 376.020 783.400 383.900 1533.320 ;
        RECT 386.100 1527.205 405.620 1533.320 ;
        RECT 407.820 1527.205 415.220 1552.545 ;
        RECT 417.420 1543.880 461.740 1552.570 ;
        RECT 463.940 1543.880 471.820 2293.800 ;
        RECT 474.020 1543.880 549.660 2293.800 ;
        RECT 551.860 1543.880 559.740 2293.800 ;
        RECT 561.940 2287.205 595.620 2293.800 ;
        RECT 597.820 2287.205 605.220 2330.070 ;
        RECT 607.420 2293.800 785.620 2330.070 ;
        RECT 607.420 2287.205 638.140 2293.800 ;
        RECT 561.940 1552.570 638.140 2287.205 ;
        RECT 561.940 1543.880 595.620 1552.570 ;
        RECT 417.420 1533.320 595.620 1543.880 ;
        RECT 417.420 1527.205 461.740 1533.320 ;
        RECT 386.100 792.570 461.740 1527.205 ;
        RECT 386.100 792.545 415.220 792.570 ;
        RECT 386.100 783.400 405.620 792.545 ;
        RECT 227.420 772.840 405.620 783.400 ;
        RECT 227.420 767.230 285.900 772.840 ;
        RECT 210.260 30.020 285.900 767.230 ;
        RECT 210.260 22.920 215.620 30.020 ;
        RECT 37.420 15.080 215.620 22.920 ;
        RECT 217.820 15.080 225.220 30.020 ;
        RECT 227.420 22.920 285.900 30.020 ;
        RECT 288.100 22.920 295.980 772.840 ;
        RECT 298.180 22.920 373.820 772.840 ;
        RECT 376.020 22.920 383.900 772.840 ;
        RECT 386.100 767.205 405.620 772.840 ;
        RECT 407.820 767.205 415.220 792.545 ;
        RECT 417.420 783.400 461.740 792.570 ;
        RECT 463.940 783.400 471.820 1533.320 ;
        RECT 474.020 783.400 549.660 1533.320 ;
        RECT 551.860 783.400 559.740 1533.320 ;
        RECT 561.940 1527.205 595.620 1533.320 ;
        RECT 597.820 1527.205 605.220 1552.570 ;
        RECT 607.420 1543.880 638.140 1552.570 ;
        RECT 640.340 1543.880 648.220 2293.800 ;
        RECT 650.420 1543.880 726.060 2293.800 ;
        RECT 728.260 1543.880 736.140 2293.800 ;
        RECT 738.340 2287.230 785.620 2293.800 ;
        RECT 787.820 2287.230 795.220 2330.070 ;
        RECT 797.420 2293.800 975.620 2330.070 ;
        RECT 797.420 2287.230 813.980 2293.800 ;
        RECT 738.340 1552.570 813.980 2287.230 ;
        RECT 738.340 1543.880 785.620 1552.570 ;
        RECT 607.420 1533.320 785.620 1543.880 ;
        RECT 607.420 1527.205 638.140 1533.320 ;
        RECT 561.940 792.570 638.140 1527.205 ;
        RECT 561.940 783.400 595.620 792.570 ;
        RECT 417.420 772.840 595.620 783.400 ;
        RECT 417.420 767.205 461.740 772.840 ;
        RECT 386.100 32.570 461.740 767.205 ;
        RECT 386.100 32.545 415.220 32.570 ;
        RECT 386.100 22.920 405.620 32.545 ;
        RECT 227.420 15.080 405.620 22.920 ;
        RECT 407.820 15.080 415.220 32.545 ;
        RECT 417.420 22.920 461.740 32.570 ;
        RECT 463.940 22.920 471.820 772.840 ;
        RECT 474.020 22.920 549.660 772.840 ;
        RECT 551.860 22.920 559.740 772.840 ;
        RECT 561.940 767.205 595.620 772.840 ;
        RECT 597.820 767.205 605.220 792.570 ;
        RECT 607.420 783.400 638.140 792.570 ;
        RECT 640.340 783.400 648.220 1533.320 ;
        RECT 650.420 783.400 726.060 1533.320 ;
        RECT 728.260 783.400 736.140 1533.320 ;
        RECT 738.340 1527.230 785.620 1533.320 ;
        RECT 787.820 1527.230 795.220 1552.570 ;
        RECT 797.420 1543.880 813.980 1552.570 ;
        RECT 816.180 1543.880 824.060 2293.800 ;
        RECT 826.260 1543.880 901.900 2293.800 ;
        RECT 904.100 1543.880 911.980 2293.800 ;
        RECT 914.180 2287.205 975.620 2293.800 ;
        RECT 977.820 2287.205 985.220 2330.070 ;
        RECT 914.180 1552.545 985.220 2287.205 ;
        RECT 914.180 1543.880 975.620 1552.545 ;
        RECT 797.420 1533.320 975.620 1543.880 ;
        RECT 797.420 1527.230 813.980 1533.320 ;
        RECT 738.340 792.570 813.980 1527.230 ;
        RECT 738.340 783.400 785.620 792.570 ;
        RECT 607.420 772.840 785.620 783.400 ;
        RECT 607.420 767.205 638.140 772.840 ;
        RECT 561.940 32.570 638.140 767.205 ;
        RECT 561.940 22.920 595.620 32.570 ;
        RECT 417.420 15.080 595.620 22.920 ;
        RECT 597.820 15.080 605.220 32.570 ;
        RECT 607.420 22.920 638.140 32.570 ;
        RECT 640.340 22.920 648.220 772.840 ;
        RECT 650.420 22.920 726.060 772.840 ;
        RECT 728.260 22.920 736.140 772.840 ;
        RECT 738.340 767.230 785.620 772.840 ;
        RECT 787.820 767.230 795.220 792.570 ;
        RECT 797.420 783.400 813.980 792.570 ;
        RECT 816.180 783.400 824.060 1533.320 ;
        RECT 826.260 783.400 901.900 1533.320 ;
        RECT 904.100 783.400 911.980 1533.320 ;
        RECT 914.180 1527.205 975.620 1533.320 ;
        RECT 977.820 1527.205 985.220 1552.545 ;
        RECT 914.180 792.545 985.220 1527.205 ;
        RECT 914.180 783.400 975.620 792.545 ;
        RECT 797.420 772.840 975.620 783.400 ;
        RECT 797.420 767.230 813.980 772.840 ;
        RECT 738.340 32.570 813.980 767.230 ;
        RECT 738.340 22.920 785.620 32.570 ;
        RECT 607.420 15.080 785.620 22.920 ;
        RECT 787.820 15.080 795.220 32.570 ;
        RECT 797.420 22.920 813.980 32.570 ;
        RECT 816.180 22.920 824.060 772.840 ;
        RECT 826.260 22.920 901.900 772.840 ;
        RECT 904.100 22.920 911.980 772.840 ;
        RECT 914.180 767.205 975.620 772.840 ;
        RECT 977.820 767.205 985.220 792.545 ;
        RECT 914.180 32.545 985.220 767.205 ;
        RECT 914.180 22.920 975.620 32.545 ;
        RECT 797.420 15.080 975.620 22.920 ;
        RECT 977.820 15.080 985.220 32.545 ;
        RECT 987.420 2293.800 1165.620 2330.070 ;
        RECT 987.420 1543.880 989.820 2293.800 ;
        RECT 992.020 1543.880 999.900 2293.800 ;
        RECT 1002.100 1543.880 1077.740 2293.800 ;
        RECT 1079.940 1543.880 1087.820 2293.800 ;
        RECT 1090.020 1543.880 1165.620 2293.800 ;
        RECT 987.420 1533.320 1165.620 1543.880 ;
        RECT 987.420 783.400 989.820 1533.320 ;
        RECT 992.020 783.400 999.900 1533.320 ;
        RECT 1002.100 783.400 1077.740 1533.320 ;
        RECT 1079.940 783.400 1087.820 1533.320 ;
        RECT 1090.020 783.400 1165.620 1533.320 ;
        RECT 987.420 772.840 1165.620 783.400 ;
        RECT 987.420 22.920 989.820 772.840 ;
        RECT 992.020 22.920 999.900 772.840 ;
        RECT 1002.100 22.920 1077.740 772.840 ;
        RECT 1079.940 22.920 1087.820 772.840 ;
        RECT 1090.020 22.920 1165.620 772.840 ;
        RECT 987.420 15.080 1165.620 22.920 ;
        RECT 1167.820 15.080 1175.220 2330.070 ;
        RECT 1177.420 2293.800 1355.620 2330.070 ;
        RECT 1177.420 1543.880 1254.140 2293.800 ;
        RECT 1256.340 1543.880 1264.220 2293.800 ;
        RECT 1266.420 2289.880 1355.620 2293.800 ;
        RECT 1266.420 1543.880 1347.100 2289.880 ;
        RECT 1349.300 1543.880 1355.620 2289.880 ;
        RECT 1177.420 1533.320 1355.620 1543.880 ;
        RECT 1177.420 783.400 1254.140 1533.320 ;
        RECT 1256.340 783.400 1264.220 1533.320 ;
        RECT 1266.420 1529.400 1355.620 1533.320 ;
        RECT 1266.420 783.400 1347.100 1529.400 ;
        RECT 1349.300 783.400 1355.620 1529.400 ;
        RECT 1177.420 772.840 1355.620 783.400 ;
        RECT 1177.420 22.920 1254.140 772.840 ;
        RECT 1256.340 22.920 1264.220 772.840 ;
        RECT 1266.420 768.920 1355.620 772.840 ;
        RECT 1266.420 22.920 1347.100 768.920 ;
        RECT 1349.300 22.920 1355.620 768.920 ;
        RECT 1177.420 15.080 1355.620 22.920 ;
        RECT 1357.820 2287.230 1365.220 2330.070 ;
        RECT 1367.420 2293.800 1545.620 2330.070 ;
        RECT 1367.420 2287.230 1429.980 2293.800 ;
        RECT 1357.820 1550.020 1429.980 2287.230 ;
        RECT 1357.820 1527.230 1365.220 1550.020 ;
        RECT 1367.420 1543.880 1429.980 1550.020 ;
        RECT 1432.180 1543.880 1440.060 2293.800 ;
        RECT 1442.260 1543.880 1517.900 2293.800 ;
        RECT 1520.100 1543.880 1527.980 2293.800 ;
        RECT 1530.180 2287.230 1545.620 2293.800 ;
        RECT 1547.820 2287.230 1555.220 2330.070 ;
        RECT 1530.180 2287.205 1555.220 2287.230 ;
        RECT 1557.420 2293.800 1735.620 2330.070 ;
        RECT 1557.420 2287.205 1605.820 2293.800 ;
        RECT 1530.180 1552.570 1605.820 2287.205 ;
        RECT 1530.180 1550.020 1555.220 1552.570 ;
        RECT 1530.180 1543.880 1545.620 1550.020 ;
        RECT 1367.420 1533.320 1545.620 1543.880 ;
        RECT 1367.420 1527.230 1429.980 1533.320 ;
        RECT 1357.820 790.020 1429.980 1527.230 ;
        RECT 1357.820 767.230 1365.220 790.020 ;
        RECT 1367.420 783.400 1429.980 790.020 ;
        RECT 1432.180 783.400 1440.060 1533.320 ;
        RECT 1442.260 783.400 1517.900 1533.320 ;
        RECT 1520.100 783.400 1527.980 1533.320 ;
        RECT 1530.180 1527.230 1545.620 1533.320 ;
        RECT 1547.820 1527.230 1555.220 1550.020 ;
        RECT 1530.180 1527.205 1555.220 1527.230 ;
        RECT 1557.420 1543.880 1605.820 1552.570 ;
        RECT 1608.020 1543.880 1615.900 2293.800 ;
        RECT 1618.100 1543.880 1693.740 2293.800 ;
        RECT 1695.940 1543.880 1703.820 2293.800 ;
        RECT 1706.020 2287.205 1735.620 2293.800 ;
        RECT 1737.820 2287.205 1745.220 2330.070 ;
        RECT 1747.420 2293.800 1925.620 2330.070 ;
        RECT 1747.420 2287.205 1781.660 2293.800 ;
        RECT 1706.020 1552.570 1781.660 2287.205 ;
        RECT 1706.020 1543.880 1735.620 1552.570 ;
        RECT 1557.420 1533.320 1735.620 1543.880 ;
        RECT 1557.420 1527.205 1605.820 1533.320 ;
        RECT 1530.180 792.570 1605.820 1527.205 ;
        RECT 1530.180 790.020 1555.220 792.570 ;
        RECT 1530.180 783.400 1545.620 790.020 ;
        RECT 1367.420 772.840 1545.620 783.400 ;
        RECT 1367.420 767.230 1429.980 772.840 ;
        RECT 1357.820 30.020 1429.980 767.230 ;
        RECT 1357.820 15.080 1365.220 30.020 ;
        RECT 1367.420 22.920 1429.980 30.020 ;
        RECT 1432.180 22.920 1440.060 772.840 ;
        RECT 1442.260 22.920 1517.900 772.840 ;
        RECT 1520.100 22.920 1527.980 772.840 ;
        RECT 1530.180 767.230 1545.620 772.840 ;
        RECT 1547.820 767.230 1555.220 790.020 ;
        RECT 1530.180 767.205 1555.220 767.230 ;
        RECT 1557.420 783.400 1605.820 792.570 ;
        RECT 1608.020 783.400 1615.900 1533.320 ;
        RECT 1618.100 783.400 1693.740 1533.320 ;
        RECT 1695.940 783.400 1703.820 1533.320 ;
        RECT 1706.020 1527.205 1735.620 1533.320 ;
        RECT 1737.820 1527.205 1745.220 1552.570 ;
        RECT 1747.420 1543.880 1781.660 1552.570 ;
        RECT 1783.860 1543.880 1791.740 2293.800 ;
        RECT 1793.940 1543.880 1870.140 2293.800 ;
        RECT 1872.340 1543.880 1880.220 2293.800 ;
        RECT 1882.420 2287.205 1925.620 2293.800 ;
        RECT 1927.820 2287.230 1935.220 2330.070 ;
        RECT 1937.420 2293.800 2115.620 2330.070 ;
        RECT 1937.420 2287.230 1958.060 2293.800 ;
        RECT 1927.820 2287.205 1958.060 2287.230 ;
        RECT 1882.420 1552.570 1958.060 2287.205 ;
        RECT 1882.420 1543.880 1925.620 1552.570 ;
        RECT 1747.420 1533.320 1925.620 1543.880 ;
        RECT 1747.420 1527.205 1781.660 1533.320 ;
        RECT 1706.020 792.570 1781.660 1527.205 ;
        RECT 1706.020 783.400 1735.620 792.570 ;
        RECT 1557.420 772.840 1735.620 783.400 ;
        RECT 1557.420 767.205 1605.820 772.840 ;
        RECT 1530.180 32.570 1605.820 767.205 ;
        RECT 1530.180 30.020 1555.220 32.570 ;
        RECT 1530.180 22.920 1545.620 30.020 ;
        RECT 1367.420 15.080 1545.620 22.920 ;
        RECT 1547.820 15.080 1555.220 30.020 ;
        RECT 1557.420 22.920 1605.820 32.570 ;
        RECT 1608.020 22.920 1615.900 772.840 ;
        RECT 1618.100 22.920 1693.740 772.840 ;
        RECT 1695.940 22.920 1703.820 772.840 ;
        RECT 1706.020 767.205 1735.620 772.840 ;
        RECT 1737.820 767.205 1745.220 792.570 ;
        RECT 1747.420 783.400 1781.660 792.570 ;
        RECT 1783.860 783.400 1791.740 1533.320 ;
        RECT 1793.940 783.400 1870.140 1533.320 ;
        RECT 1872.340 783.400 1880.220 1533.320 ;
        RECT 1882.420 1527.205 1925.620 1533.320 ;
        RECT 1927.820 1527.230 1935.220 1552.570 ;
        RECT 1937.420 1543.880 1958.060 1552.570 ;
        RECT 1960.260 1543.880 1968.140 2293.800 ;
        RECT 1970.340 1543.880 2045.980 2293.800 ;
        RECT 2048.180 1543.880 2056.060 2293.800 ;
        RECT 2058.260 2287.230 2115.620 2293.800 ;
        RECT 2117.820 2287.815 2125.220 2330.070 ;
        RECT 2127.420 2293.800 2147.460 2330.070 ;
        RECT 2127.420 2287.815 2143.420 2293.800 ;
        RECT 2117.820 2287.230 2143.420 2287.815 ;
        RECT 2058.260 1552.545 2143.420 2287.230 ;
        RECT 2058.260 1543.880 2115.620 1552.545 ;
        RECT 1937.420 1533.320 2115.620 1543.880 ;
        RECT 1937.420 1527.230 1958.060 1533.320 ;
        RECT 1927.820 1527.205 1958.060 1527.230 ;
        RECT 1882.420 792.570 1958.060 1527.205 ;
        RECT 1882.420 783.400 1925.620 792.570 ;
        RECT 1747.420 772.840 1925.620 783.400 ;
        RECT 1747.420 767.205 1781.660 772.840 ;
        RECT 1706.020 32.570 1781.660 767.205 ;
        RECT 1706.020 22.920 1735.620 32.570 ;
        RECT 1557.420 15.080 1735.620 22.920 ;
        RECT 1737.820 15.080 1745.220 32.570 ;
        RECT 1747.420 22.920 1781.660 32.570 ;
        RECT 1783.860 22.920 1791.740 772.840 ;
        RECT 1793.940 22.920 1870.140 772.840 ;
        RECT 1872.340 22.920 1880.220 772.840 ;
        RECT 1882.420 767.205 1925.620 772.840 ;
        RECT 1927.820 767.230 1935.220 792.570 ;
        RECT 1937.420 783.400 1958.060 792.570 ;
        RECT 1960.260 783.400 1968.140 1533.320 ;
        RECT 1970.340 783.400 2045.980 1533.320 ;
        RECT 2048.180 783.400 2056.060 1533.320 ;
        RECT 2058.260 1527.230 2115.620 1533.320 ;
        RECT 2117.820 1550.810 2143.420 1552.545 ;
        RECT 2117.820 1527.815 2125.220 1550.810 ;
        RECT 2127.420 1543.880 2143.420 1550.810 ;
        RECT 2145.620 1543.880 2147.460 2293.800 ;
        RECT 2127.420 1533.320 2147.460 1543.880 ;
        RECT 2127.420 1527.815 2143.420 1533.320 ;
        RECT 2117.820 1527.230 2143.420 1527.815 ;
        RECT 2058.260 792.545 2143.420 1527.230 ;
        RECT 2058.260 783.400 2115.620 792.545 ;
        RECT 1937.420 772.840 2115.620 783.400 ;
        RECT 1937.420 767.230 1958.060 772.840 ;
        RECT 1927.820 767.205 1958.060 767.230 ;
        RECT 1882.420 32.570 1958.060 767.205 ;
        RECT 1882.420 22.920 1925.620 32.570 ;
        RECT 1747.420 15.080 1925.620 22.920 ;
        RECT 1927.820 15.080 1935.220 32.570 ;
        RECT 1937.420 22.920 1958.060 32.570 ;
        RECT 1960.260 22.920 1968.140 772.840 ;
        RECT 1970.340 22.920 2045.980 772.840 ;
        RECT 2048.180 22.920 2056.060 772.840 ;
        RECT 2058.260 767.230 2115.620 772.840 ;
        RECT 2117.820 790.810 2143.420 792.545 ;
        RECT 2117.820 767.815 2125.220 790.810 ;
        RECT 2127.420 783.400 2143.420 790.810 ;
        RECT 2145.620 783.400 2147.460 1533.320 ;
        RECT 2127.420 772.840 2147.460 783.400 ;
        RECT 2127.420 767.815 2143.420 772.840 ;
        RECT 2117.820 767.230 2143.420 767.815 ;
        RECT 2058.260 32.545 2143.420 767.230 ;
        RECT 2058.260 22.920 2115.620 32.545 ;
        RECT 1937.420 15.080 2115.620 22.920 ;
        RECT 2117.820 30.810 2143.420 32.545 ;
        RECT 2117.820 15.080 2125.220 30.810 ;
        RECT 2127.420 22.920 2143.420 30.810 ;
        RECT 2145.620 22.920 2147.460 772.840 ;
        RECT 2127.420 15.080 2147.460 22.920 ;
        RECT 16.940 1.210 2147.460 15.080 ;
      LAYER Metal5 ;
        RECT 10 0 2165 34.5 ;
        RECT 10 49.5 2165 79.5 ;
        RECT 10 94.5 2165 124.5 ;
        RECT 10 139.5 2165 169.5 ;
        RECT 10 184.5 2165 214.5 ;
        RECT 10 229.5 2165 259.5 ;
        RECT 10 274.5 2165 304.5 ;
        RECT 10 319.5 2165 349.5 ;
        RECT 10 364.5 2165 394.5 ;
        RECT 10 409.5 2165 439.5 ;
        RECT 10 454.5 2165 484.5 ;
        RECT 10 499.5 2165 529.5 ;
        RECT 10 544.5 2165 574.5 ;
        RECT 10 589.5 2165 619.5 ;
        RECT 10 634.5 2165 664.5 ;
        RECT 10 679.5 2165 709.5 ;
        RECT 10 724.5 2165 754.5 ;
        RECT 10 769.5 2165 799.5 ;
        RECT 10 814.5 2165 844.5 ;
        RECT 10 859.5 2165 889.5 ;
        RECT 10 904.5 2165 934.5 ;
        RECT 10 949.5 2165 979.5 ;
        RECT 10 994.5 2165 1024.5 ;
        RECT 10 1039.5 2165 1069.5 ;
        RECT 10 1084.5 2165 1114.5 ;
        RECT 10 1129.5 2165 1159.5 ;
        RECT 10 1174.5 2165 1204.5 ;
        RECT 10 1219.5 2165 1249.5 ;
        RECT 10 1264.5 2165 1294.5 ;
        RECT 10 1309.5 2165 1339.5 ;
        RECT 10 1354.5 2165 1384.5 ;
        RECT 10 1399.5 2165 1429.5 ;
        RECT 10 1444.5 2165 1474.5 ;
        RECT 10 1489.5 2165 1519.5 ;
        RECT 10 1534.5 2165 1564.5 ;
        RECT 10 1579.5 2165 1609.5 ;
        RECT 10 1624.5 2165 1654.5 ;
        RECT 10 1669.5 2165 1699.5 ;
        RECT 10 1714.5 2165 1744.5 ;
        RECT 10 1759.5 2165 1789.5 ;
        RECT 10 1804.5 2165 1834.5 ;
        RECT 10 1849.5 2165 1879.5 ;
        RECT 10 1894.5 2165 1924.5 ;
        RECT 10 1939.5 2165 1969.5 ;
        RECT 10 1984.5 2165 2014.5 ;
        RECT 10 2029.5 2165 2059.5 ;
        RECT 10 2074.5 2165 2104.5 ;
        RECT 10 2119.5 2165 2149.5 ;
        RECT 10 2164.5 2165 2194.5 ;
        RECT 10 2209.5 2165 2239.5 ;
        RECT 10 2254.5 2165 2284.5 ;
        RECT 10 2299.5 2165 2329.5 ;
  END
END efuse_ctrl
END LIBRARY

