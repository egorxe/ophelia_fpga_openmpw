VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2980.200 BY 2980.200 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 35.560 2985.000 36.680 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2017.960 2985.000 2019.080 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2216.200 2985.000 2217.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2414.440 2985.000 2415.560 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2612.680 2985.000 2613.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2810.920 2985.000 2812.040 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2923.480 2977.800 2924.600 2985.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2592.520 2977.800 2593.640 2985.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2261.560 2977.800 2262.680 2985.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1930.600 2977.800 1931.720 2985.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1599.640 2977.800 1600.760 2985.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 233.800 2985.000 234.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.680 2977.800 1269.800 2985.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.720 2977.800 938.840 2985.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 606.760 2977.800 607.880 2985.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 2977.800 276.920 2985.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2935.800 2.400 2936.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2724.120 2.400 2725.240 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2512.440 2.400 2513.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2300.760 2.400 2301.880 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2089.080 2.400 2090.200 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1877.400 2.400 1878.520 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 432.040 2985.000 433.160 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1665.720 2.400 1666.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1454.040 2.400 1455.160 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1242.360 2.400 1243.480 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1030.680 2.400 1031.800 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 819.000 2.400 820.120 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 607.320 2.400 608.440 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 395.640 2.400 396.760 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 183.960 2.400 185.080 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 630.280 2985.000 631.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 828.520 2985.000 829.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1026.760 2985.000 1027.880 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1225.000 2985.000 1226.120 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1423.240 2985.000 1424.360 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1621.480 2985.000 1622.600 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1819.720 2985.000 1820.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 167.720 2985.000 168.840 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2150.120 2985.000 2151.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2348.360 2985.000 2349.480 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2546.600 2985.000 2547.720 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2744.840 2985.000 2745.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2943.080 2985.000 2944.200 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2702.840 2977.800 2703.960 2985.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2371.880 2977.800 2373.000 2985.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2040.920 2977.800 2042.040 2985.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1709.960 2977.800 1711.080 2985.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1379.000 2977.800 1380.120 2985.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 365.960 2985.000 367.080 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.040 2977.800 1049.160 2985.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 717.080 2977.800 718.200 2985.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.120 2977.800 387.240 2985.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 2977.800 56.280 2985.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2794.680 2.400 2795.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2583.000 2.400 2584.120 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2371.320 2.400 2372.440 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2159.640 2.400 2160.760 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1947.960 2.400 1949.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1736.280 2.400 1737.400 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 564.200 2985.000 565.320 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1524.600 2.400 1525.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1312.920 2.400 1314.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1101.240 2.400 1102.360 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 889.560 2.400 890.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 677.880 2.400 679.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 466.200 2.400 467.320 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 254.520 2.400 255.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 42.840 2.400 43.960 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 762.440 2985.000 763.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 960.680 2985.000 961.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1158.920 2985.000 1160.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1357.160 2985.000 1358.280 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1555.400 2985.000 1556.520 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1753.640 2985.000 1754.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1951.880 2985.000 1953.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 101.640 2985.000 102.760 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2084.040 2985.000 2085.160 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2282.280 2985.000 2283.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2480.520 2985.000 2481.640 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2678.760 2985.000 2679.880 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2877.000 2985.000 2878.120 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2813.160 2977.800 2814.280 2985.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2482.200 2977.800 2483.320 2985.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2151.240 2977.800 2152.360 2985.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1820.280 2977.800 1821.400 2985.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1489.320 2977.800 1490.440 2985.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 299.880 2985.000 301.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1158.360 2977.800 1159.480 2985.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 827.400 2977.800 828.520 2985.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.440 2977.800 497.560 2985.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.480 2977.800 166.600 2985.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2865.240 2.400 2866.360 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2653.560 2.400 2654.680 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2441.880 2.400 2443.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2230.200 2.400 2231.320 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2018.520 2.400 2019.640 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1806.840 2.400 1807.960 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 498.120 2985.000 499.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1595.160 2.400 1596.280 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1383.480 2.400 1384.600 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1171.800 2.400 1172.920 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 960.120 2.400 961.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 748.440 2.400 749.560 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 536.760 2.400 537.880 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 325.080 2.400 326.200 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 113.400 2.400 114.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 696.360 2985.000 697.480 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 894.600 2985.000 895.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1092.840 2985.000 1093.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1291.080 2985.000 1292.200 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1489.320 2985.000 1490.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1687.560 2985.000 1688.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1885.800 2985.000 1886.920 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.960 -4.800 1067.080 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1351.560 -4.800 1352.680 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1380.120 -4.800 1381.240 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1408.680 -4.800 1409.800 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1437.240 -4.800 1438.360 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1465.800 -4.800 1466.920 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1494.360 -4.800 1495.480 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1522.920 -4.800 1524.040 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1551.480 -4.800 1552.600 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1580.040 -4.800 1581.160 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1608.600 -4.800 1609.720 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1094.520 -4.800 1095.640 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1637.160 -4.800 1638.280 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1665.720 -4.800 1666.840 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1694.280 -4.800 1695.400 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1722.840 -4.800 1723.960 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1751.400 -4.800 1752.520 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1779.960 -4.800 1781.080 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.520 -4.800 1809.640 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1837.080 -4.800 1838.200 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1865.640 -4.800 1866.760 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1894.200 -4.800 1895.320 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1123.080 -4.800 1124.200 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1922.760 -4.800 1923.880 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1951.320 -4.800 1952.440 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1979.880 -4.800 1981.000 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2008.440 -4.800 2009.560 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2037.000 -4.800 2038.120 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2065.560 -4.800 2066.680 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2094.120 -4.800 2095.240 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2122.680 -4.800 2123.800 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2151.240 -4.800 2152.360 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2179.800 -4.800 2180.920 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1151.640 -4.800 1152.760 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2208.360 -4.800 2209.480 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2236.920 -4.800 2238.040 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2265.480 -4.800 2266.600 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2294.040 -4.800 2295.160 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2322.600 -4.800 2323.720 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2351.160 -4.800 2352.280 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2379.720 -4.800 2380.840 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2408.280 -4.800 2409.400 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2436.840 -4.800 2437.960 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2465.400 -4.800 2466.520 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1180.200 -4.800 1181.320 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2493.960 -4.800 2495.080 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2522.520 -4.800 2523.640 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2551.080 -4.800 2552.200 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2579.640 -4.800 2580.760 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2608.200 -4.800 2609.320 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2636.760 -4.800 2637.880 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2665.320 -4.800 2666.440 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2693.880 -4.800 2695.000 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2722.440 -4.800 2723.560 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2751.000 -4.800 2752.120 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1208.760 -4.800 1209.880 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2779.560 -4.800 2780.680 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2808.120 -4.800 2809.240 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2836.680 -4.800 2837.800 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2865.240 -4.800 2866.360 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1237.320 -4.800 1238.440 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1265.880 -4.800 1267.000 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1294.440 -4.800 1295.560 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1323.000 -4.800 1324.120 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1075.480 -4.800 1076.600 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1361.080 -4.800 1362.200 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1389.640 -4.800 1390.760 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1418.200 -4.800 1419.320 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1446.760 -4.800 1447.880 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1475.320 -4.800 1476.440 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1503.880 -4.800 1505.000 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1532.440 -4.800 1533.560 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1561.000 -4.800 1562.120 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1589.560 -4.800 1590.680 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1618.120 -4.800 1619.240 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1104.040 -4.800 1105.160 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1646.680 -4.800 1647.800 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1675.240 -4.800 1676.360 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1703.800 -4.800 1704.920 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1732.360 -4.800 1733.480 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1760.920 -4.800 1762.040 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1789.480 -4.800 1790.600 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.040 -4.800 1819.160 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1846.600 -4.800 1847.720 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1875.160 -4.800 1876.280 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1903.720 -4.800 1904.840 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.600 -4.800 1133.720 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1932.280 -4.800 1933.400 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1960.840 -4.800 1961.960 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1989.400 -4.800 1990.520 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2017.960 -4.800 2019.080 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2046.520 -4.800 2047.640 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2075.080 -4.800 2076.200 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2103.640 -4.800 2104.760 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2132.200 -4.800 2133.320 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2160.760 -4.800 2161.880 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.320 -4.800 2190.440 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1161.160 -4.800 1162.280 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2217.880 -4.800 2219.000 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2246.440 -4.800 2247.560 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2275.000 -4.800 2276.120 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2303.560 -4.800 2304.680 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2332.120 -4.800 2333.240 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2360.680 -4.800 2361.800 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2389.240 -4.800 2390.360 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2417.800 -4.800 2418.920 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2446.360 -4.800 2447.480 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2474.920 -4.800 2476.040 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1189.720 -4.800 1190.840 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2503.480 -4.800 2504.600 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2532.040 -4.800 2533.160 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2560.600 -4.800 2561.720 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2589.160 -4.800 2590.280 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2617.720 -4.800 2618.840 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2646.280 -4.800 2647.400 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2674.840 -4.800 2675.960 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2703.400 -4.800 2704.520 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2731.960 -4.800 2733.080 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2760.520 -4.800 2761.640 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1218.280 -4.800 1219.400 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2789.080 -4.800 2790.200 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2817.640 -4.800 2818.760 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2846.200 -4.800 2847.320 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2874.760 -4.800 2875.880 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1246.840 -4.800 1247.960 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.400 -4.800 1276.520 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1303.960 -4.800 1305.080 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.520 -4.800 1333.640 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1085.000 -4.800 1086.120 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1370.600 -4.800 1371.720 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1399.160 -4.800 1400.280 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1427.720 -4.800 1428.840 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1456.280 -4.800 1457.400 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.840 -4.800 1485.960 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1513.400 -4.800 1514.520 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1541.960 -4.800 1543.080 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1570.520 -4.800 1571.640 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1599.080 -4.800 1600.200 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1627.640 -4.800 1628.760 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1113.560 -4.800 1114.680 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1656.200 -4.800 1657.320 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1684.760 -4.800 1685.880 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1713.320 -4.800 1714.440 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1741.880 -4.800 1743.000 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1770.440 -4.800 1771.560 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1799.000 -4.800 1800.120 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1827.560 -4.800 1828.680 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1856.120 -4.800 1857.240 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1884.680 -4.800 1885.800 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1913.240 -4.800 1914.360 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1142.120 -4.800 1143.240 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1941.800 -4.800 1942.920 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.360 -4.800 1971.480 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1998.920 -4.800 2000.040 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2027.480 -4.800 2028.600 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2056.040 -4.800 2057.160 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2084.600 -4.800 2085.720 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2113.160 -4.800 2114.280 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2141.720 -4.800 2142.840 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2170.280 -4.800 2171.400 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2198.840 -4.800 2199.960 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1170.680 -4.800 1171.800 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2227.400 -4.800 2228.520 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2255.960 -4.800 2257.080 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2284.520 -4.800 2285.640 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2313.080 -4.800 2314.200 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2341.640 -4.800 2342.760 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.200 -4.800 2371.320 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2398.760 -4.800 2399.880 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.320 -4.800 2428.440 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2455.880 -4.800 2457.000 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2484.440 -4.800 2485.560 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1199.240 -4.800 1200.360 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2513.000 -4.800 2514.120 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2541.560 -4.800 2542.680 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2570.120 -4.800 2571.240 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2598.680 -4.800 2599.800 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2627.240 -4.800 2628.360 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2655.800 -4.800 2656.920 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2684.360 -4.800 2685.480 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2712.920 -4.800 2714.040 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2741.480 -4.800 2742.600 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2770.040 -4.800 2771.160 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1227.800 -4.800 1228.920 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2798.600 -4.800 2799.720 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2827.160 -4.800 2828.280 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2855.720 -4.800 2856.840 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2884.280 -4.800 2885.400 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1256.360 -4.800 1257.480 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1284.920 -4.800 1286.040 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1313.480 -4.800 1314.600 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1342.040 -4.800 1343.160 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2893.800 -4.800 2894.920 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2903.320 -4.800 2904.440 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2912.840 -4.800 2913.960 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2922.360 -4.800 2923.480 2.400 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -4.780 -3.420 -1.680 2986.540 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 -3.420 2985.100 -0.320 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 2983.440 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2982.000 -3.420 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.770 -8.220 18.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 -8.220 128.870 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 390.950 128.870 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 810.950 128.870 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 1230.950 128.870 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 1650.950 128.870 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 2070.950 128.870 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 2490.950 128.870 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 125.770 2910.950 128.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 -8.220 238.870 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 390.950 238.870 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 810.950 238.870 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 1230.950 238.870 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 1650.950 238.870 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 2070.950 238.870 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 2490.950 238.870 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.770 2910.950 238.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 345.770 -8.220 348.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 -8.220 458.870 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 390.950 458.870 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 810.950 458.870 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 1230.950 458.870 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 1650.950 458.870 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 2070.950 458.870 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 2490.950 458.870 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 455.770 2910.950 458.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 -8.220 568.870 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 390.950 568.870 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 810.950 568.870 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 1230.950 568.870 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 1650.950 568.870 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 2070.950 568.870 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 2490.950 568.870 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.770 2910.950 568.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 675.770 -8.220 678.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.770 -8.220 788.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.770 2864.815 788.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 895.770 -8.220 898.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 895.770 2864.815 898.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1005.770 -8.220 1008.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1005.770 2864.815 1008.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1115.770 -8.220 1118.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1115.770 2880.080 1118.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1225.770 -8.220 1228.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1225.770 2864.815 1228.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1335.770 -8.220 1338.870 571.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1335.770 2919.280 1338.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1445.770 -8.220 1448.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1445.770 2864.815 1448.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.770 -8.220 1558.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.770 2880.080 1558.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1665.770 -8.220 1668.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1665.770 2864.815 1668.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1775.770 -8.220 1778.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1775.770 2864.815 1778.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1885.770 -8.220 1888.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1885.770 2864.815 1888.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1995.770 -8.220 1998.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1995.770 2880.080 1998.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2105.770 -8.220 2108.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2105.770 2864.815 2108.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2215.770 -8.220 2218.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2215.770 2864.815 2218.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2325.770 -8.220 2328.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2325.770 2864.815 2328.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2435.770 -8.220 2438.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2435.770 2880.080 2438.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2545.770 -8.220 2548.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2545.770 2864.815 2548.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2655.770 -8.220 2658.870 571.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2655.770 2919.280 2658.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2765.770 -8.220 2768.870 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2765.770 2864.815 2768.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2875.770 -8.220 2878.870 599.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2875.770 2880.080 2878.870 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 17.130 2989.900 20.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 107.130 2989.900 110.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 197.130 2989.900 200.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 287.130 2989.900 290.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 377.130 2989.900 380.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 467.130 2989.900 470.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 557.130 736.240 560.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 647.130 2989.900 650.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 737.130 2989.900 740.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 827.130 2989.900 830.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 917.130 2989.900 920.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1007.130 2989.900 1010.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1097.130 2989.900 1100.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1187.130 2989.900 1190.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1277.130 2989.900 1280.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1367.130 2989.900 1370.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1457.130 2989.900 1460.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1547.130 2989.900 1550.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1637.130 2989.900 1640.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1727.130 2989.900 1730.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1817.130 2989.900 1820.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1907.130 2989.900 1910.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1997.130 2989.900 2000.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2087.130 2989.900 2090.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2177.130 2989.900 2180.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2267.130 2989.900 2270.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2357.130 2989.900 2360.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2447.130 2989.900 2450.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2537.130 2989.900 2540.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2627.130 2989.900 2630.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2717.130 2989.900 2720.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2807.130 2989.900 2810.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2897.130 2989.900 2900.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2902.160 557.130 2989.900 560.230 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2934.250 544.580 2937.350 2948.140 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -9.580 -8.220 -6.480 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 -8.220 2989.900 -5.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2988.240 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.800 -8.220 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.870 -8.220 31.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 -8.220 141.970 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 390.950 141.970 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 810.950 141.970 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 1230.950 141.970 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 1650.950 141.970 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 2070.950 141.970 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 2490.950 141.970 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.870 2910.950 141.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 -8.220 251.970 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 390.950 251.970 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 810.950 251.970 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 1230.950 251.970 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 1650.950 251.970 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 2070.950 251.970 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 2490.950 251.970 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.870 2910.950 251.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.870 -8.220 361.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 -8.220 471.970 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 390.950 471.970 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 810.950 471.970 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 1230.950 471.970 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 1650.950 471.970 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 2070.950 471.970 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 2490.950 471.970 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 468.870 2910.950 471.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 -8.220 581.970 80.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 390.950 581.970 500.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 810.950 581.970 920.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 1230.950 581.970 1340.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 1650.950 581.970 1760.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 2070.950 581.970 2180.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 2490.950 581.970 2600.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.870 2910.950 581.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.870 -8.220 691.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 798.870 -8.220 801.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 798.870 2864.815 801.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 908.870 -8.220 911.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 908.870 2864.815 911.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1018.870 -8.220 1021.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1018.870 2880.080 1021.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1128.870 -8.220 1131.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1128.870 2864.815 1131.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1238.870 -8.220 1241.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1238.870 2864.815 1241.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1348.870 -8.220 1351.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1348.870 2864.815 1351.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1458.870 -8.220 1461.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1458.870 2880.080 1461.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.870 -8.220 1571.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.870 2864.815 1571.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1678.870 -8.220 1681.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1678.870 2864.815 1681.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.870 -8.220 1791.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.870 2864.815 1791.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1898.870 -8.220 1901.970 571.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1898.870 2919.280 1901.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2008.870 -8.220 2011.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2008.870 2864.815 2011.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2118.870 -8.220 2121.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2118.870 2864.815 2121.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2228.870 -8.220 2231.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2228.870 2864.815 2231.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2338.870 -8.220 2341.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2338.870 2880.080 2341.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.870 -8.220 2451.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.870 2864.815 2451.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2558.870 -8.220 2561.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2558.870 2864.815 2561.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2668.870 -8.220 2671.970 571.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2668.870 2919.280 2671.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2778.870 -8.220 2781.970 574.430 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2778.870 2880.080 2781.970 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2888.870 -8.220 2891.970 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 62.130 2989.900 65.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 152.130 2989.900 155.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 242.130 2989.900 245.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 332.130 2989.900 335.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 422.130 2989.900 425.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 512.130 2989.900 515.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 602.130 2989.900 605.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 692.130 2989.900 695.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 782.130 2989.900 785.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 872.130 2989.900 875.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 962.130 2989.900 965.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1052.130 2989.900 1055.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1142.130 2989.900 1145.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1232.130 2989.900 1235.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1322.130 2989.900 1325.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1412.130 2989.900 1415.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1502.130 2989.900 1505.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1592.130 2989.900 1595.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1682.130 2989.900 1685.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1772.130 2989.900 1775.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1862.130 2989.900 1865.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1952.130 2989.900 1955.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2042.130 2989.900 2045.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2132.130 2989.900 2135.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2222.130 2989.900 2225.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2312.130 2989.900 2315.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2402.130 2989.900 2405.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2492.130 2989.900 2495.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2582.130 2989.900 2585.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2672.130 2989.900 2675.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2762.130 2989.900 2765.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2852.130 2989.900 2855.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2942.130 2989.900 2945.230 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2947.690 544.580 2950.790 2948.140 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 -4.800 57.960 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.360 -4.800 67.480 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.880 -4.800 77.000 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 -4.800 115.080 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.640 -4.800 438.760 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.200 -4.800 467.320 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.760 -4.800 495.880 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.320 -4.800 524.440 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.880 -4.800 553.000 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.440 -4.800 581.560 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.000 -4.800 610.120 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 637.560 -4.800 638.680 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 666.120 -4.800 667.240 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 694.680 -4.800 695.800 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.040 -4.800 153.160 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.240 -4.800 724.360 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.800 -4.800 752.920 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 780.360 -4.800 781.480 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.920 -4.800 810.040 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.480 -4.800 838.600 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.040 -4.800 867.160 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.600 -4.800 895.720 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 923.160 -4.800 924.280 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 951.720 -4.800 952.840 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 980.280 -4.800 981.400 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.120 -4.800 191.240 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1008.840 -4.800 1009.960 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.400 -4.800 1038.520 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 -4.800 229.320 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.280 -4.800 267.400 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 -4.800 295.960 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.400 -4.800 324.520 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 -4.800 353.080 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.520 -4.800 381.640 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.080 -4.800 410.200 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.400 -4.800 86.520 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 -4.800 124.600 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.160 -4.800 448.280 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 475.720 -4.800 476.840 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.280 -4.800 505.400 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.840 -4.800 533.960 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.400 -4.800 562.520 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 589.960 -4.800 591.080 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.520 -4.800 619.640 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.080 -4.800 648.200 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.640 -4.800 676.760 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 704.200 -4.800 705.320 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 -4.800 162.680 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.760 -4.800 733.880 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 761.320 -4.800 762.440 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.880 -4.800 791.000 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 818.440 -4.800 819.560 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.000 -4.800 848.120 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.560 -4.800 876.680 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 904.120 -4.800 905.240 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 932.680 -4.800 933.800 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 961.240 -4.800 962.360 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 989.800 -4.800 990.920 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.640 -4.800 200.760 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.360 -4.800 1019.480 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1046.920 -4.800 1048.040 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 -4.800 238.840 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 -4.800 276.920 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.360 -4.800 305.480 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.920 -4.800 334.040 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.480 -4.800 362.600 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.040 -4.800 391.160 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.600 -4.800 419.720 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.000 -4.800 134.120 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.680 -4.800 457.800 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 485.240 -4.800 486.360 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.800 -4.800 514.920 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.360 -4.800 543.480 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.920 -4.800 572.040 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.480 -4.800 600.600 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.040 -4.800 629.160 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 656.600 -4.800 657.720 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.160 -4.800 686.280 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 713.720 -4.800 714.840 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.080 -4.800 172.200 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.280 -4.800 743.400 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.840 -4.800 771.960 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.400 -4.800 800.520 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 827.960 -4.800 829.080 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.520 -4.800 857.640 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 885.080 -4.800 886.200 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.640 -4.800 914.760 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 942.200 -4.800 943.320 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 970.760 -4.800 971.880 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 999.320 -4.800 1000.440 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.160 -4.800 210.280 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1027.880 -4.800 1029.000 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.440 -4.800 1057.560 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.240 -4.800 248.360 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.320 -4.800 286.440 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.880 -4.800 315.000 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.440 -4.800 343.560 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 -4.800 372.120 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.560 -4.800 400.680 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.120 -4.800 429.240 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.520 -4.800 143.640 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 -4.800 181.720 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.680 -4.800 219.800 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 -4.800 257.880 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.920 -4.800 96.040 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 -4.800 105.560 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 8.490 14.710 2968.000 2968.410 ;
      LAYER Metal2 ;
        RECT 0.140 2977.500 54.860 2979.670 ;
        RECT 56.580 2977.500 165.180 2979.670 ;
        RECT 166.900 2977.500 275.500 2979.670 ;
        RECT 277.220 2977.500 385.820 2979.670 ;
        RECT 387.540 2977.500 496.140 2979.670 ;
        RECT 497.860 2977.500 606.460 2979.670 ;
        RECT 608.180 2977.500 716.780 2979.670 ;
        RECT 718.500 2977.500 827.100 2979.670 ;
        RECT 828.820 2977.500 937.420 2979.670 ;
        RECT 939.140 2977.500 1047.740 2979.670 ;
        RECT 1049.460 2977.500 1158.060 2979.670 ;
        RECT 1159.780 2977.500 1268.380 2979.670 ;
        RECT 1270.100 2977.500 1378.700 2979.670 ;
        RECT 1380.420 2977.500 1489.020 2979.670 ;
        RECT 1490.740 2977.500 1599.340 2979.670 ;
        RECT 1601.060 2977.500 1709.660 2979.670 ;
        RECT 1711.380 2977.500 1819.980 2979.670 ;
        RECT 1821.700 2977.500 1930.300 2979.670 ;
        RECT 1932.020 2977.500 2040.620 2979.670 ;
        RECT 2042.340 2977.500 2150.940 2979.670 ;
        RECT 2152.660 2977.500 2261.260 2979.670 ;
        RECT 2262.980 2977.500 2371.580 2979.670 ;
        RECT 2373.300 2977.500 2481.900 2979.670 ;
        RECT 2483.620 2977.500 2592.220 2979.670 ;
        RECT 2593.940 2977.500 2702.540 2979.670 ;
        RECT 2704.260 2977.500 2812.860 2979.670 ;
        RECT 2814.580 2977.500 2923.180 2979.670 ;
        RECT 2924.900 2977.500 2965.620 2979.670 ;
        RECT 0.140 2.700 2965.620 2977.500 ;
        RECT 0.140 1.770 56.540 2.700 ;
        RECT 58.260 1.770 66.060 2.700 ;
        RECT 67.780 1.770 75.580 2.700 ;
        RECT 77.300 1.770 85.100 2.700 ;
        RECT 86.820 1.770 94.620 2.700 ;
        RECT 96.340 1.770 104.140 2.700 ;
        RECT 105.860 1.770 113.660 2.700 ;
        RECT 115.380 1.770 123.180 2.700 ;
        RECT 124.900 1.770 132.700 2.700 ;
        RECT 134.420 1.770 142.220 2.700 ;
        RECT 143.940 1.770 151.740 2.700 ;
        RECT 153.460 1.770 161.260 2.700 ;
        RECT 162.980 1.770 170.780 2.700 ;
        RECT 172.500 1.770 180.300 2.700 ;
        RECT 182.020 1.770 189.820 2.700 ;
        RECT 191.540 1.770 199.340 2.700 ;
        RECT 201.060 1.770 208.860 2.700 ;
        RECT 210.580 1.770 218.380 2.700 ;
        RECT 220.100 1.770 227.900 2.700 ;
        RECT 229.620 1.770 237.420 2.700 ;
        RECT 239.140 1.770 246.940 2.700 ;
        RECT 248.660 1.770 256.460 2.700 ;
        RECT 258.180 1.770 265.980 2.700 ;
        RECT 267.700 1.770 275.500 2.700 ;
        RECT 277.220 1.770 285.020 2.700 ;
        RECT 286.740 1.770 294.540 2.700 ;
        RECT 296.260 1.770 304.060 2.700 ;
        RECT 305.780 1.770 313.580 2.700 ;
        RECT 315.300 1.770 323.100 2.700 ;
        RECT 324.820 1.770 332.620 2.700 ;
        RECT 334.340 1.770 342.140 2.700 ;
        RECT 343.860 1.770 351.660 2.700 ;
        RECT 353.380 1.770 361.180 2.700 ;
        RECT 362.900 1.770 370.700 2.700 ;
        RECT 372.420 1.770 380.220 2.700 ;
        RECT 381.940 1.770 389.740 2.700 ;
        RECT 391.460 1.770 399.260 2.700 ;
        RECT 400.980 1.770 408.780 2.700 ;
        RECT 410.500 1.770 418.300 2.700 ;
        RECT 420.020 1.770 427.820 2.700 ;
        RECT 429.540 1.770 437.340 2.700 ;
        RECT 439.060 1.770 446.860 2.700 ;
        RECT 448.580 1.770 456.380 2.700 ;
        RECT 458.100 1.770 465.900 2.700 ;
        RECT 467.620 1.770 475.420 2.700 ;
        RECT 477.140 1.770 484.940 2.700 ;
        RECT 486.660 1.770 494.460 2.700 ;
        RECT 496.180 1.770 503.980 2.700 ;
        RECT 505.700 1.770 513.500 2.700 ;
        RECT 515.220 1.770 523.020 2.700 ;
        RECT 524.740 1.770 532.540 2.700 ;
        RECT 534.260 1.770 542.060 2.700 ;
        RECT 543.780 1.770 551.580 2.700 ;
        RECT 553.300 1.770 561.100 2.700 ;
        RECT 562.820 1.770 570.620 2.700 ;
        RECT 572.340 1.770 580.140 2.700 ;
        RECT 581.860 1.770 589.660 2.700 ;
        RECT 591.380 1.770 599.180 2.700 ;
        RECT 600.900 1.770 608.700 2.700 ;
        RECT 610.420 1.770 618.220 2.700 ;
        RECT 619.940 1.770 627.740 2.700 ;
        RECT 629.460 1.770 637.260 2.700 ;
        RECT 638.980 1.770 646.780 2.700 ;
        RECT 648.500 1.770 656.300 2.700 ;
        RECT 658.020 1.770 665.820 2.700 ;
        RECT 667.540 1.770 675.340 2.700 ;
        RECT 677.060 1.770 684.860 2.700 ;
        RECT 686.580 1.770 694.380 2.700 ;
        RECT 696.100 1.770 703.900 2.700 ;
        RECT 705.620 1.770 713.420 2.700 ;
        RECT 715.140 1.770 722.940 2.700 ;
        RECT 724.660 1.770 732.460 2.700 ;
        RECT 734.180 1.770 741.980 2.700 ;
        RECT 743.700 1.770 751.500 2.700 ;
        RECT 753.220 1.770 761.020 2.700 ;
        RECT 762.740 1.770 770.540 2.700 ;
        RECT 772.260 1.770 780.060 2.700 ;
        RECT 781.780 1.770 789.580 2.700 ;
        RECT 791.300 1.770 799.100 2.700 ;
        RECT 800.820 1.770 808.620 2.700 ;
        RECT 810.340 1.770 818.140 2.700 ;
        RECT 819.860 1.770 827.660 2.700 ;
        RECT 829.380 1.770 837.180 2.700 ;
        RECT 838.900 1.770 846.700 2.700 ;
        RECT 848.420 1.770 856.220 2.700 ;
        RECT 857.940 1.770 865.740 2.700 ;
        RECT 867.460 1.770 875.260 2.700 ;
        RECT 876.980 1.770 884.780 2.700 ;
        RECT 886.500 1.770 894.300 2.700 ;
        RECT 896.020 1.770 903.820 2.700 ;
        RECT 905.540 1.770 913.340 2.700 ;
        RECT 915.060 1.770 922.860 2.700 ;
        RECT 924.580 1.770 932.380 2.700 ;
        RECT 934.100 1.770 941.900 2.700 ;
        RECT 943.620 1.770 951.420 2.700 ;
        RECT 953.140 1.770 960.940 2.700 ;
        RECT 962.660 1.770 970.460 2.700 ;
        RECT 972.180 1.770 979.980 2.700 ;
        RECT 981.700 1.770 989.500 2.700 ;
        RECT 991.220 1.770 999.020 2.700 ;
        RECT 1000.740 1.770 1008.540 2.700 ;
        RECT 1010.260 1.770 1018.060 2.700 ;
        RECT 1019.780 1.770 1027.580 2.700 ;
        RECT 1029.300 1.770 1037.100 2.700 ;
        RECT 1038.820 1.770 1046.620 2.700 ;
        RECT 1048.340 1.770 1056.140 2.700 ;
        RECT 1057.860 1.770 1065.660 2.700 ;
        RECT 1067.380 1.770 1075.180 2.700 ;
        RECT 1076.900 1.770 1084.700 2.700 ;
        RECT 1086.420 1.770 1094.220 2.700 ;
        RECT 1095.940 1.770 1103.740 2.700 ;
        RECT 1105.460 1.770 1113.260 2.700 ;
        RECT 1114.980 1.770 1122.780 2.700 ;
        RECT 1124.500 1.770 1132.300 2.700 ;
        RECT 1134.020 1.770 1141.820 2.700 ;
        RECT 1143.540 1.770 1151.340 2.700 ;
        RECT 1153.060 1.770 1160.860 2.700 ;
        RECT 1162.580 1.770 1170.380 2.700 ;
        RECT 1172.100 1.770 1179.900 2.700 ;
        RECT 1181.620 1.770 1189.420 2.700 ;
        RECT 1191.140 1.770 1198.940 2.700 ;
        RECT 1200.660 1.770 1208.460 2.700 ;
        RECT 1210.180 1.770 1217.980 2.700 ;
        RECT 1219.700 1.770 1227.500 2.700 ;
        RECT 1229.220 1.770 1237.020 2.700 ;
        RECT 1238.740 1.770 1246.540 2.700 ;
        RECT 1248.260 1.770 1256.060 2.700 ;
        RECT 1257.780 1.770 1265.580 2.700 ;
        RECT 1267.300 1.770 1275.100 2.700 ;
        RECT 1276.820 1.770 1284.620 2.700 ;
        RECT 1286.340 1.770 1294.140 2.700 ;
        RECT 1295.860 1.770 1303.660 2.700 ;
        RECT 1305.380 1.770 1313.180 2.700 ;
        RECT 1314.900 1.770 1322.700 2.700 ;
        RECT 1324.420 1.770 1332.220 2.700 ;
        RECT 1333.940 1.770 1341.740 2.700 ;
        RECT 1343.460 1.770 1351.260 2.700 ;
        RECT 1352.980 1.770 1360.780 2.700 ;
        RECT 1362.500 1.770 1370.300 2.700 ;
        RECT 1372.020 1.770 1379.820 2.700 ;
        RECT 1381.540 1.770 1389.340 2.700 ;
        RECT 1391.060 1.770 1398.860 2.700 ;
        RECT 1400.580 1.770 1408.380 2.700 ;
        RECT 1410.100 1.770 1417.900 2.700 ;
        RECT 1419.620 1.770 1427.420 2.700 ;
        RECT 1429.140 1.770 1436.940 2.700 ;
        RECT 1438.660 1.770 1446.460 2.700 ;
        RECT 1448.180 1.770 1455.980 2.700 ;
        RECT 1457.700 1.770 1465.500 2.700 ;
        RECT 1467.220 1.770 1475.020 2.700 ;
        RECT 1476.740 1.770 1484.540 2.700 ;
        RECT 1486.260 1.770 1494.060 2.700 ;
        RECT 1495.780 1.770 1503.580 2.700 ;
        RECT 1505.300 1.770 1513.100 2.700 ;
        RECT 1514.820 1.770 1522.620 2.700 ;
        RECT 1524.340 1.770 1532.140 2.700 ;
        RECT 1533.860 1.770 1541.660 2.700 ;
        RECT 1543.380 1.770 1551.180 2.700 ;
        RECT 1552.900 1.770 1560.700 2.700 ;
        RECT 1562.420 1.770 1570.220 2.700 ;
        RECT 1571.940 1.770 1579.740 2.700 ;
        RECT 1581.460 1.770 1589.260 2.700 ;
        RECT 1590.980 1.770 1598.780 2.700 ;
        RECT 1600.500 1.770 1608.300 2.700 ;
        RECT 1610.020 1.770 1617.820 2.700 ;
        RECT 1619.540 1.770 1627.340 2.700 ;
        RECT 1629.060 1.770 1636.860 2.700 ;
        RECT 1638.580 1.770 1646.380 2.700 ;
        RECT 1648.100 1.770 1655.900 2.700 ;
        RECT 1657.620 1.770 1665.420 2.700 ;
        RECT 1667.140 1.770 1674.940 2.700 ;
        RECT 1676.660 1.770 1684.460 2.700 ;
        RECT 1686.180 1.770 1693.980 2.700 ;
        RECT 1695.700 1.770 1703.500 2.700 ;
        RECT 1705.220 1.770 1713.020 2.700 ;
        RECT 1714.740 1.770 1722.540 2.700 ;
        RECT 1724.260 1.770 1732.060 2.700 ;
        RECT 1733.780 1.770 1741.580 2.700 ;
        RECT 1743.300 1.770 1751.100 2.700 ;
        RECT 1752.820 1.770 1760.620 2.700 ;
        RECT 1762.340 1.770 1770.140 2.700 ;
        RECT 1771.860 1.770 1779.660 2.700 ;
        RECT 1781.380 1.770 1789.180 2.700 ;
        RECT 1790.900 1.770 1798.700 2.700 ;
        RECT 1800.420 1.770 1808.220 2.700 ;
        RECT 1809.940 1.770 1817.740 2.700 ;
        RECT 1819.460 1.770 1827.260 2.700 ;
        RECT 1828.980 1.770 1836.780 2.700 ;
        RECT 1838.500 1.770 1846.300 2.700 ;
        RECT 1848.020 1.770 1855.820 2.700 ;
        RECT 1857.540 1.770 1865.340 2.700 ;
        RECT 1867.060 1.770 1874.860 2.700 ;
        RECT 1876.580 1.770 1884.380 2.700 ;
        RECT 1886.100 1.770 1893.900 2.700 ;
        RECT 1895.620 1.770 1903.420 2.700 ;
        RECT 1905.140 1.770 1912.940 2.700 ;
        RECT 1914.660 1.770 1922.460 2.700 ;
        RECT 1924.180 1.770 1931.980 2.700 ;
        RECT 1933.700 1.770 1941.500 2.700 ;
        RECT 1943.220 1.770 1951.020 2.700 ;
        RECT 1952.740 1.770 1960.540 2.700 ;
        RECT 1962.260 1.770 1970.060 2.700 ;
        RECT 1971.780 1.770 1979.580 2.700 ;
        RECT 1981.300 1.770 1989.100 2.700 ;
        RECT 1990.820 1.770 1998.620 2.700 ;
        RECT 2000.340 1.770 2008.140 2.700 ;
        RECT 2009.860 1.770 2017.660 2.700 ;
        RECT 2019.380 1.770 2027.180 2.700 ;
        RECT 2028.900 1.770 2036.700 2.700 ;
        RECT 2038.420 1.770 2046.220 2.700 ;
        RECT 2047.940 1.770 2055.740 2.700 ;
        RECT 2057.460 1.770 2065.260 2.700 ;
        RECT 2066.980 1.770 2074.780 2.700 ;
        RECT 2076.500 1.770 2084.300 2.700 ;
        RECT 2086.020 1.770 2093.820 2.700 ;
        RECT 2095.540 1.770 2103.340 2.700 ;
        RECT 2105.060 1.770 2112.860 2.700 ;
        RECT 2114.580 1.770 2122.380 2.700 ;
        RECT 2124.100 1.770 2131.900 2.700 ;
        RECT 2133.620 1.770 2141.420 2.700 ;
        RECT 2143.140 1.770 2150.940 2.700 ;
        RECT 2152.660 1.770 2160.460 2.700 ;
        RECT 2162.180 1.770 2169.980 2.700 ;
        RECT 2171.700 1.770 2179.500 2.700 ;
        RECT 2181.220 1.770 2189.020 2.700 ;
        RECT 2190.740 1.770 2198.540 2.700 ;
        RECT 2200.260 1.770 2208.060 2.700 ;
        RECT 2209.780 1.770 2217.580 2.700 ;
        RECT 2219.300 1.770 2227.100 2.700 ;
        RECT 2228.820 1.770 2236.620 2.700 ;
        RECT 2238.340 1.770 2246.140 2.700 ;
        RECT 2247.860 1.770 2255.660 2.700 ;
        RECT 2257.380 1.770 2265.180 2.700 ;
        RECT 2266.900 1.770 2274.700 2.700 ;
        RECT 2276.420 1.770 2284.220 2.700 ;
        RECT 2285.940 1.770 2293.740 2.700 ;
        RECT 2295.460 1.770 2303.260 2.700 ;
        RECT 2304.980 1.770 2312.780 2.700 ;
        RECT 2314.500 1.770 2322.300 2.700 ;
        RECT 2324.020 1.770 2331.820 2.700 ;
        RECT 2333.540 1.770 2341.340 2.700 ;
        RECT 2343.060 1.770 2350.860 2.700 ;
        RECT 2352.580 1.770 2360.380 2.700 ;
        RECT 2362.100 1.770 2369.900 2.700 ;
        RECT 2371.620 1.770 2379.420 2.700 ;
        RECT 2381.140 1.770 2388.940 2.700 ;
        RECT 2390.660 1.770 2398.460 2.700 ;
        RECT 2400.180 1.770 2407.980 2.700 ;
        RECT 2409.700 1.770 2417.500 2.700 ;
        RECT 2419.220 1.770 2427.020 2.700 ;
        RECT 2428.740 1.770 2436.540 2.700 ;
        RECT 2438.260 1.770 2446.060 2.700 ;
        RECT 2447.780 1.770 2455.580 2.700 ;
        RECT 2457.300 1.770 2465.100 2.700 ;
        RECT 2466.820 1.770 2474.620 2.700 ;
        RECT 2476.340 1.770 2484.140 2.700 ;
        RECT 2485.860 1.770 2493.660 2.700 ;
        RECT 2495.380 1.770 2503.180 2.700 ;
        RECT 2504.900 1.770 2512.700 2.700 ;
        RECT 2514.420 1.770 2522.220 2.700 ;
        RECT 2523.940 1.770 2531.740 2.700 ;
        RECT 2533.460 1.770 2541.260 2.700 ;
        RECT 2542.980 1.770 2550.780 2.700 ;
        RECT 2552.500 1.770 2560.300 2.700 ;
        RECT 2562.020 1.770 2569.820 2.700 ;
        RECT 2571.540 1.770 2579.340 2.700 ;
        RECT 2581.060 1.770 2588.860 2.700 ;
        RECT 2590.580 1.770 2598.380 2.700 ;
        RECT 2600.100 1.770 2607.900 2.700 ;
        RECT 2609.620 1.770 2617.420 2.700 ;
        RECT 2619.140 1.770 2626.940 2.700 ;
        RECT 2628.660 1.770 2636.460 2.700 ;
        RECT 2638.180 1.770 2645.980 2.700 ;
        RECT 2647.700 1.770 2655.500 2.700 ;
        RECT 2657.220 1.770 2665.020 2.700 ;
        RECT 2666.740 1.770 2674.540 2.700 ;
        RECT 2676.260 1.770 2684.060 2.700 ;
        RECT 2685.780 1.770 2693.580 2.700 ;
        RECT 2695.300 1.770 2703.100 2.700 ;
        RECT 2704.820 1.770 2712.620 2.700 ;
        RECT 2714.340 1.770 2722.140 2.700 ;
        RECT 2723.860 1.770 2731.660 2.700 ;
        RECT 2733.380 1.770 2741.180 2.700 ;
        RECT 2742.900 1.770 2750.700 2.700 ;
        RECT 2752.420 1.770 2760.220 2.700 ;
        RECT 2761.940 1.770 2769.740 2.700 ;
        RECT 2771.460 1.770 2779.260 2.700 ;
        RECT 2780.980 1.770 2788.780 2.700 ;
        RECT 2790.500 1.770 2798.300 2.700 ;
        RECT 2800.020 1.770 2807.820 2.700 ;
        RECT 2809.540 1.770 2817.340 2.700 ;
        RECT 2819.060 1.770 2826.860 2.700 ;
        RECT 2828.580 1.770 2836.380 2.700 ;
        RECT 2838.100 1.770 2845.900 2.700 ;
        RECT 2847.620 1.770 2855.420 2.700 ;
        RECT 2857.140 1.770 2864.940 2.700 ;
        RECT 2866.660 1.770 2874.460 2.700 ;
        RECT 2876.180 1.770 2883.980 2.700 ;
        RECT 2885.700 1.770 2893.500 2.700 ;
        RECT 2895.220 1.770 2903.020 2.700 ;
        RECT 2904.740 1.770 2912.540 2.700 ;
        RECT 2914.260 1.770 2922.060 2.700 ;
        RECT 2923.780 1.770 2965.620 2.700 ;
      LAYER Metal3 ;
        RECT 0.090 2944.500 2978.360 2979.620 ;
        RECT 0.090 2942.780 2977.500 2944.500 ;
        RECT 0.090 2937.220 2978.360 2942.780 ;
        RECT 2.700 2935.500 2978.360 2937.220 ;
        RECT 0.090 2878.420 2978.360 2935.500 ;
        RECT 0.090 2876.700 2977.500 2878.420 ;
        RECT 0.090 2866.660 2978.360 2876.700 ;
        RECT 2.700 2864.940 2978.360 2866.660 ;
        RECT 0.090 2812.340 2978.360 2864.940 ;
        RECT 0.090 2810.620 2977.500 2812.340 ;
        RECT 0.090 2796.100 2978.360 2810.620 ;
        RECT 2.700 2794.380 2978.360 2796.100 ;
        RECT 0.090 2746.260 2978.360 2794.380 ;
        RECT 0.090 2744.540 2977.500 2746.260 ;
        RECT 0.090 2725.540 2978.360 2744.540 ;
        RECT 2.700 2723.820 2978.360 2725.540 ;
        RECT 0.090 2680.180 2978.360 2723.820 ;
        RECT 0.090 2678.460 2977.500 2680.180 ;
        RECT 0.090 2654.980 2978.360 2678.460 ;
        RECT 2.700 2653.260 2978.360 2654.980 ;
        RECT 0.090 2614.100 2978.360 2653.260 ;
        RECT 0.090 2612.380 2977.500 2614.100 ;
        RECT 0.090 2584.420 2978.360 2612.380 ;
        RECT 2.700 2582.700 2978.360 2584.420 ;
        RECT 0.090 2548.020 2978.360 2582.700 ;
        RECT 0.090 2546.300 2977.500 2548.020 ;
        RECT 0.090 2513.860 2978.360 2546.300 ;
        RECT 2.700 2512.140 2978.360 2513.860 ;
        RECT 0.090 2481.940 2978.360 2512.140 ;
        RECT 0.090 2480.220 2977.500 2481.940 ;
        RECT 0.090 2443.300 2978.360 2480.220 ;
        RECT 2.700 2441.580 2978.360 2443.300 ;
        RECT 0.090 2415.860 2978.360 2441.580 ;
        RECT 0.090 2414.140 2977.500 2415.860 ;
        RECT 0.090 2372.740 2978.360 2414.140 ;
        RECT 2.700 2371.020 2978.360 2372.740 ;
        RECT 0.090 2349.780 2978.360 2371.020 ;
        RECT 0.090 2348.060 2977.500 2349.780 ;
        RECT 0.090 2302.180 2978.360 2348.060 ;
        RECT 2.700 2300.460 2978.360 2302.180 ;
        RECT 0.090 2283.700 2978.360 2300.460 ;
        RECT 0.090 2281.980 2977.500 2283.700 ;
        RECT 0.090 2231.620 2978.360 2281.980 ;
        RECT 2.700 2229.900 2978.360 2231.620 ;
        RECT 0.090 2217.620 2978.360 2229.900 ;
        RECT 0.090 2215.900 2977.500 2217.620 ;
        RECT 0.090 2161.060 2978.360 2215.900 ;
        RECT 2.700 2159.340 2978.360 2161.060 ;
        RECT 0.090 2151.540 2978.360 2159.340 ;
        RECT 0.090 2149.820 2977.500 2151.540 ;
        RECT 0.090 2090.500 2978.360 2149.820 ;
        RECT 2.700 2088.780 2978.360 2090.500 ;
        RECT 0.090 2085.460 2978.360 2088.780 ;
        RECT 0.090 2083.740 2977.500 2085.460 ;
        RECT 0.090 2019.940 2978.360 2083.740 ;
        RECT 2.700 2019.380 2978.360 2019.940 ;
        RECT 2.700 2018.220 2977.500 2019.380 ;
        RECT 0.090 2017.660 2977.500 2018.220 ;
        RECT 0.090 1953.300 2978.360 2017.660 ;
        RECT 0.090 1951.580 2977.500 1953.300 ;
        RECT 0.090 1949.380 2978.360 1951.580 ;
        RECT 2.700 1947.660 2978.360 1949.380 ;
        RECT 0.090 1887.220 2978.360 1947.660 ;
        RECT 0.090 1885.500 2977.500 1887.220 ;
        RECT 0.090 1878.820 2978.360 1885.500 ;
        RECT 2.700 1877.100 2978.360 1878.820 ;
        RECT 0.090 1821.140 2978.360 1877.100 ;
        RECT 0.090 1819.420 2977.500 1821.140 ;
        RECT 0.090 1808.260 2978.360 1819.420 ;
        RECT 2.700 1806.540 2978.360 1808.260 ;
        RECT 0.090 1755.060 2978.360 1806.540 ;
        RECT 0.090 1753.340 2977.500 1755.060 ;
        RECT 0.090 1737.700 2978.360 1753.340 ;
        RECT 2.700 1735.980 2978.360 1737.700 ;
        RECT 0.090 1688.980 2978.360 1735.980 ;
        RECT 0.090 1687.260 2977.500 1688.980 ;
        RECT 0.090 1667.140 2978.360 1687.260 ;
        RECT 2.700 1665.420 2978.360 1667.140 ;
        RECT 0.090 1622.900 2978.360 1665.420 ;
        RECT 0.090 1621.180 2977.500 1622.900 ;
        RECT 0.090 1596.580 2978.360 1621.180 ;
        RECT 2.700 1594.860 2978.360 1596.580 ;
        RECT 0.090 1556.820 2978.360 1594.860 ;
        RECT 0.090 1555.100 2977.500 1556.820 ;
        RECT 0.090 1526.020 2978.360 1555.100 ;
        RECT 2.700 1524.300 2978.360 1526.020 ;
        RECT 0.090 1490.740 2978.360 1524.300 ;
        RECT 0.090 1489.020 2977.500 1490.740 ;
        RECT 0.090 1455.460 2978.360 1489.020 ;
        RECT 2.700 1453.740 2978.360 1455.460 ;
        RECT 0.090 1424.660 2978.360 1453.740 ;
        RECT 0.090 1422.940 2977.500 1424.660 ;
        RECT 0.090 1384.900 2978.360 1422.940 ;
        RECT 2.700 1383.180 2978.360 1384.900 ;
        RECT 0.090 1358.580 2978.360 1383.180 ;
        RECT 0.090 1356.860 2977.500 1358.580 ;
        RECT 0.090 1314.340 2978.360 1356.860 ;
        RECT 2.700 1312.620 2978.360 1314.340 ;
        RECT 0.090 1292.500 2978.360 1312.620 ;
        RECT 0.090 1290.780 2977.500 1292.500 ;
        RECT 0.090 1243.780 2978.360 1290.780 ;
        RECT 2.700 1242.060 2978.360 1243.780 ;
        RECT 0.090 1226.420 2978.360 1242.060 ;
        RECT 0.090 1224.700 2977.500 1226.420 ;
        RECT 0.090 1173.220 2978.360 1224.700 ;
        RECT 2.700 1171.500 2978.360 1173.220 ;
        RECT 0.090 1160.340 2978.360 1171.500 ;
        RECT 0.090 1158.620 2977.500 1160.340 ;
        RECT 0.090 1102.660 2978.360 1158.620 ;
        RECT 2.700 1100.940 2978.360 1102.660 ;
        RECT 0.090 1094.260 2978.360 1100.940 ;
        RECT 0.090 1092.540 2977.500 1094.260 ;
        RECT 0.090 1032.100 2978.360 1092.540 ;
        RECT 2.700 1030.380 2978.360 1032.100 ;
        RECT 0.090 1028.180 2978.360 1030.380 ;
        RECT 0.090 1026.460 2977.500 1028.180 ;
        RECT 0.090 962.100 2978.360 1026.460 ;
        RECT 0.090 961.540 2977.500 962.100 ;
        RECT 2.700 960.380 2977.500 961.540 ;
        RECT 2.700 959.820 2978.360 960.380 ;
        RECT 0.090 896.020 2978.360 959.820 ;
        RECT 0.090 894.300 2977.500 896.020 ;
        RECT 0.090 890.980 2978.360 894.300 ;
        RECT 2.700 889.260 2978.360 890.980 ;
        RECT 0.090 829.940 2978.360 889.260 ;
        RECT 0.090 828.220 2977.500 829.940 ;
        RECT 0.090 820.420 2978.360 828.220 ;
        RECT 2.700 818.700 2978.360 820.420 ;
        RECT 0.090 763.860 2978.360 818.700 ;
        RECT 0.090 762.140 2977.500 763.860 ;
        RECT 0.090 749.860 2978.360 762.140 ;
        RECT 2.700 748.140 2978.360 749.860 ;
        RECT 0.090 697.780 2978.360 748.140 ;
        RECT 0.090 696.060 2977.500 697.780 ;
        RECT 0.090 679.300 2978.360 696.060 ;
        RECT 2.700 677.580 2978.360 679.300 ;
        RECT 0.090 631.700 2978.360 677.580 ;
        RECT 0.090 629.980 2977.500 631.700 ;
        RECT 0.090 608.740 2978.360 629.980 ;
        RECT 2.700 607.020 2978.360 608.740 ;
        RECT 0.090 565.620 2978.360 607.020 ;
        RECT 0.090 563.900 2977.500 565.620 ;
        RECT 0.090 538.180 2978.360 563.900 ;
        RECT 2.700 536.460 2978.360 538.180 ;
        RECT 0.090 499.540 2978.360 536.460 ;
        RECT 0.090 497.820 2977.500 499.540 ;
        RECT 0.090 467.620 2978.360 497.820 ;
        RECT 2.700 465.900 2978.360 467.620 ;
        RECT 0.090 433.460 2978.360 465.900 ;
        RECT 0.090 431.740 2977.500 433.460 ;
        RECT 0.090 397.060 2978.360 431.740 ;
        RECT 2.700 395.340 2978.360 397.060 ;
        RECT 0.090 367.380 2978.360 395.340 ;
        RECT 0.090 365.660 2977.500 367.380 ;
        RECT 0.090 326.500 2978.360 365.660 ;
        RECT 2.700 324.780 2978.360 326.500 ;
        RECT 0.090 301.300 2978.360 324.780 ;
        RECT 0.090 299.580 2977.500 301.300 ;
        RECT 0.090 255.940 2978.360 299.580 ;
        RECT 2.700 254.220 2978.360 255.940 ;
        RECT 0.090 235.220 2978.360 254.220 ;
        RECT 0.090 233.500 2977.500 235.220 ;
        RECT 0.090 185.380 2978.360 233.500 ;
        RECT 2.700 183.660 2978.360 185.380 ;
        RECT 0.090 169.140 2978.360 183.660 ;
        RECT 0.090 167.420 2977.500 169.140 ;
        RECT 0.090 114.820 2978.360 167.420 ;
        RECT 2.700 113.100 2978.360 114.820 ;
        RECT 0.090 103.060 2978.360 113.100 ;
        RECT 0.090 101.340 2977.500 103.060 ;
        RECT 0.090 44.260 2978.360 101.340 ;
        RECT 2.700 42.540 2978.360 44.260 ;
        RECT 0.090 36.980 2978.360 42.540 ;
        RECT 0.090 35.260 2977.500 36.980 ;
        RECT 0.090 1.260 2978.360 35.260 ;
      LAYER Metal4 ;
        RECT 0.140 1.070 15.470 2976.870 ;
        RECT 19.170 1.070 28.570 2976.870 ;
        RECT 32.270 2910.650 125.470 2976.870 ;
        RECT 129.170 2910.650 138.570 2976.870 ;
        RECT 142.270 2910.650 235.470 2976.870 ;
        RECT 239.170 2910.650 248.570 2976.870 ;
        RECT 252.270 2910.650 345.470 2976.870 ;
        RECT 32.270 2601.270 345.470 2910.650 ;
        RECT 32.270 2490.650 125.470 2601.270 ;
        RECT 129.170 2490.650 138.570 2601.270 ;
        RECT 142.270 2490.650 235.470 2601.270 ;
        RECT 239.170 2490.650 248.570 2601.270 ;
        RECT 252.270 2490.650 345.470 2601.270 ;
        RECT 32.270 2181.270 345.470 2490.650 ;
        RECT 32.270 2070.650 125.470 2181.270 ;
        RECT 129.170 2070.650 138.570 2181.270 ;
        RECT 142.270 2070.650 235.470 2181.270 ;
        RECT 239.170 2070.650 248.570 2181.270 ;
        RECT 252.270 2070.650 345.470 2181.270 ;
        RECT 32.270 1761.270 345.470 2070.650 ;
        RECT 32.270 1650.650 125.470 1761.270 ;
        RECT 129.170 1650.650 138.570 1761.270 ;
        RECT 142.270 1650.650 235.470 1761.270 ;
        RECT 239.170 1650.650 248.570 1761.270 ;
        RECT 252.270 1650.650 345.470 1761.270 ;
        RECT 32.270 1341.270 345.470 1650.650 ;
        RECT 32.270 1230.650 125.470 1341.270 ;
        RECT 129.170 1230.650 138.570 1341.270 ;
        RECT 142.270 1230.650 235.470 1341.270 ;
        RECT 239.170 1230.650 248.570 1341.270 ;
        RECT 252.270 1230.650 345.470 1341.270 ;
        RECT 32.270 921.270 345.470 1230.650 ;
        RECT 32.270 810.650 125.470 921.270 ;
        RECT 129.170 810.650 138.570 921.270 ;
        RECT 142.270 810.650 235.470 921.270 ;
        RECT 239.170 810.650 248.570 921.270 ;
        RECT 252.270 810.650 345.470 921.270 ;
        RECT 32.270 501.270 345.470 810.650 ;
        RECT 32.270 390.650 125.470 501.270 ;
        RECT 129.170 390.650 138.570 501.270 ;
        RECT 142.270 390.650 235.470 501.270 ;
        RECT 239.170 390.650 248.570 501.270 ;
        RECT 252.270 390.650 345.470 501.270 ;
        RECT 32.270 81.270 345.470 390.650 ;
        RECT 32.270 1.070 125.470 81.270 ;
        RECT 129.170 1.070 138.570 81.270 ;
        RECT 142.270 1.070 235.470 81.270 ;
        RECT 239.170 1.070 248.570 81.270 ;
        RECT 252.270 1.070 345.470 81.270 ;
        RECT 349.170 1.070 358.570 2976.870 ;
        RECT 362.270 2910.650 455.470 2976.870 ;
        RECT 459.170 2910.650 468.570 2976.870 ;
        RECT 472.270 2910.650 565.470 2976.870 ;
        RECT 569.170 2910.650 578.570 2976.870 ;
        RECT 582.270 2910.650 675.470 2976.870 ;
        RECT 362.270 2601.270 675.470 2910.650 ;
        RECT 362.270 2490.650 455.470 2601.270 ;
        RECT 459.170 2490.650 468.570 2601.270 ;
        RECT 472.270 2490.650 565.470 2601.270 ;
        RECT 569.170 2490.650 578.570 2601.270 ;
        RECT 582.270 2490.650 675.470 2601.270 ;
        RECT 362.270 2181.270 675.470 2490.650 ;
        RECT 362.270 2070.650 455.470 2181.270 ;
        RECT 459.170 2070.650 468.570 2181.270 ;
        RECT 472.270 2070.650 565.470 2181.270 ;
        RECT 569.170 2070.650 578.570 2181.270 ;
        RECT 582.270 2070.650 675.470 2181.270 ;
        RECT 362.270 1761.270 675.470 2070.650 ;
        RECT 362.270 1650.650 455.470 1761.270 ;
        RECT 459.170 1650.650 468.570 1761.270 ;
        RECT 472.270 1650.650 565.470 1761.270 ;
        RECT 569.170 1650.650 578.570 1761.270 ;
        RECT 582.270 1650.650 675.470 1761.270 ;
        RECT 362.270 1341.270 675.470 1650.650 ;
        RECT 362.270 1230.650 455.470 1341.270 ;
        RECT 459.170 1230.650 468.570 1341.270 ;
        RECT 472.270 1230.650 565.470 1341.270 ;
        RECT 569.170 1230.650 578.570 1341.270 ;
        RECT 582.270 1230.650 675.470 1341.270 ;
        RECT 362.270 921.270 675.470 1230.650 ;
        RECT 362.270 810.650 455.470 921.270 ;
        RECT 459.170 810.650 468.570 921.270 ;
        RECT 472.270 810.650 565.470 921.270 ;
        RECT 569.170 810.650 578.570 921.270 ;
        RECT 582.270 810.650 675.470 921.270 ;
        RECT 362.270 501.270 675.470 810.650 ;
        RECT 362.270 390.650 455.470 501.270 ;
        RECT 459.170 390.650 468.570 501.270 ;
        RECT 472.270 390.650 565.470 501.270 ;
        RECT 569.170 390.650 578.570 501.270 ;
        RECT 582.270 390.650 675.470 501.270 ;
        RECT 362.270 81.270 675.470 390.650 ;
        RECT 362.270 1.070 455.470 81.270 ;
        RECT 459.170 1.070 468.570 81.270 ;
        RECT 472.270 1.070 565.470 81.270 ;
        RECT 569.170 1.070 578.570 81.270 ;
        RECT 582.270 1.070 675.470 81.270 ;
        RECT 679.170 1.070 688.570 2976.870 ;
        RECT 692.270 2864.515 785.470 2976.870 ;
        RECT 789.170 2864.515 798.570 2976.870 ;
        RECT 802.270 2864.515 895.470 2976.870 ;
        RECT 899.170 2864.515 908.570 2976.870 ;
        RECT 912.270 2864.515 1005.470 2976.870 ;
        RECT 1009.170 2879.780 1018.570 2976.870 ;
        RECT 1022.270 2879.780 1115.470 2976.870 ;
        RECT 1119.170 2879.780 1128.570 2976.870 ;
        RECT 1009.170 2864.515 1128.570 2879.780 ;
        RECT 1132.270 2864.515 1225.470 2976.870 ;
        RECT 1229.170 2864.515 1238.570 2976.870 ;
        RECT 1242.270 2918.980 1335.470 2976.870 ;
        RECT 1339.170 2918.980 1348.570 2976.870 ;
        RECT 1242.270 2864.515 1348.570 2918.980 ;
        RECT 1352.270 2864.515 1445.470 2976.870 ;
        RECT 1449.170 2879.780 1458.570 2976.870 ;
        RECT 1462.270 2879.780 1555.470 2976.870 ;
        RECT 1559.170 2879.780 1568.570 2976.870 ;
        RECT 1449.170 2864.515 1568.570 2879.780 ;
        RECT 1572.270 2864.515 1665.470 2976.870 ;
        RECT 1669.170 2864.515 1678.570 2976.870 ;
        RECT 1682.270 2864.515 1775.470 2976.870 ;
        RECT 1779.170 2864.515 1788.570 2976.870 ;
        RECT 1792.270 2864.515 1885.470 2976.870 ;
        RECT 1889.170 2918.980 1898.570 2976.870 ;
        RECT 1902.270 2918.980 1995.470 2976.870 ;
        RECT 1889.170 2879.780 1995.470 2918.980 ;
        RECT 1999.170 2879.780 2008.570 2976.870 ;
        RECT 1889.170 2864.515 2008.570 2879.780 ;
        RECT 2012.270 2864.515 2105.470 2976.870 ;
        RECT 2109.170 2864.515 2118.570 2976.870 ;
        RECT 2122.270 2864.515 2215.470 2976.870 ;
        RECT 2219.170 2864.515 2228.570 2976.870 ;
        RECT 2232.270 2864.515 2325.470 2976.870 ;
        RECT 2329.170 2879.780 2338.570 2976.870 ;
        RECT 2342.270 2879.780 2435.470 2976.870 ;
        RECT 2439.170 2879.780 2448.570 2976.870 ;
        RECT 2329.170 2864.515 2448.570 2879.780 ;
        RECT 2452.270 2864.515 2545.470 2976.870 ;
        RECT 2549.170 2864.515 2558.570 2976.870 ;
        RECT 2562.270 2918.980 2655.470 2976.870 ;
        RECT 2659.170 2918.980 2668.570 2976.870 ;
        RECT 2672.270 2918.980 2765.470 2976.870 ;
        RECT 2562.270 2864.515 2765.470 2918.980 ;
        RECT 2769.170 2879.780 2778.570 2976.870 ;
        RECT 2782.270 2879.780 2875.470 2976.870 ;
        RECT 2879.170 2879.780 2888.570 2976.870 ;
        RECT 2769.170 2864.515 2888.570 2879.780 ;
        RECT 692.270 599.540 2888.570 2864.515 ;
        RECT 692.270 574.730 2875.470 599.540 ;
        RECT 692.270 1.070 785.470 574.730 ;
        RECT 789.170 1.070 798.570 574.730 ;
        RECT 802.270 1.070 895.470 574.730 ;
        RECT 899.170 1.070 908.570 574.730 ;
        RECT 912.270 1.070 1005.470 574.730 ;
        RECT 1009.170 1.070 1018.570 574.730 ;
        RECT 1022.270 1.070 1115.470 574.730 ;
        RECT 1119.170 1.070 1128.570 574.730 ;
        RECT 1132.270 1.070 1225.470 574.730 ;
        RECT 1229.170 1.070 1238.570 574.730 ;
        RECT 1242.270 572.100 1348.570 574.730 ;
        RECT 1242.270 1.070 1335.470 572.100 ;
        RECT 1339.170 1.070 1348.570 572.100 ;
        RECT 1352.270 1.070 1445.470 574.730 ;
        RECT 1449.170 1.070 1458.570 574.730 ;
        RECT 1462.270 1.070 1555.470 574.730 ;
        RECT 1559.170 1.070 1568.570 574.730 ;
        RECT 1572.270 1.070 1665.470 574.730 ;
        RECT 1669.170 1.070 1678.570 574.730 ;
        RECT 1682.270 1.070 1775.470 574.730 ;
        RECT 1779.170 1.070 1788.570 574.730 ;
        RECT 1792.270 1.070 1885.470 574.730 ;
        RECT 1889.170 572.100 1995.470 574.730 ;
        RECT 1889.170 1.070 1898.570 572.100 ;
        RECT 1902.270 1.070 1995.470 572.100 ;
        RECT 1999.170 1.070 2008.570 574.730 ;
        RECT 2012.270 1.070 2105.470 574.730 ;
        RECT 2109.170 1.070 2118.570 574.730 ;
        RECT 2122.270 1.070 2215.470 574.730 ;
        RECT 2219.170 1.070 2228.570 574.730 ;
        RECT 2232.270 1.070 2325.470 574.730 ;
        RECT 2329.170 1.070 2338.570 574.730 ;
        RECT 2342.270 1.070 2435.470 574.730 ;
        RECT 2439.170 1.070 2448.570 574.730 ;
        RECT 2452.270 1.070 2545.470 574.730 ;
        RECT 2549.170 1.070 2558.570 574.730 ;
        RECT 2562.270 572.100 2765.470 574.730 ;
        RECT 2562.270 1.070 2655.470 572.100 ;
        RECT 2659.170 1.070 2668.570 572.100 ;
        RECT 2672.270 1.070 2765.470 572.100 ;
        RECT 2769.170 1.070 2778.570 574.730 ;
        RECT 2782.270 1.070 2875.470 574.730 ;
        RECT 2879.170 1.070 2888.570 599.540 ;
        RECT 2892.270 2948.440 2956.100 2976.870 ;
        RECT 2892.270 544.280 2933.950 2948.440 ;
        RECT 2937.650 544.280 2947.390 2948.440 ;
        RECT 2951.090 544.280 2956.100 2948.440 ;
        RECT 2892.270 1.070 2956.100 544.280 ;
      LAYER Metal5 ;
        RECT 0.060 2945.730 2956.180 2964.580 ;
        RECT 0.060 2900.730 2956.180 2941.630 ;
        RECT 0.060 2855.730 2956.180 2896.630 ;
        RECT 0.060 2810.730 2956.180 2851.630 ;
        RECT 0.060 2765.730 2956.180 2806.630 ;
        RECT 0.060 2720.730 2956.180 2761.630 ;
        RECT 0.060 2675.730 2956.180 2716.630 ;
        RECT 0.060 2630.730 2956.180 2671.630 ;
        RECT 0.060 2585.730 2956.180 2626.630 ;
        RECT 0.060 2540.730 2956.180 2581.630 ;
        RECT 0.060 2495.730 2956.180 2536.630 ;
        RECT 0.060 2450.730 2956.180 2491.630 ;
        RECT 0.060 2405.730 2956.180 2446.630 ;
        RECT 0.060 2360.730 2956.180 2401.630 ;
        RECT 0.060 2315.730 2956.180 2356.630 ;
        RECT 0.060 2270.730 2956.180 2311.630 ;
        RECT 0.060 2225.730 2956.180 2266.630 ;
        RECT 0.060 2180.730 2956.180 2221.630 ;
        RECT 0.060 2135.730 2956.180 2176.630 ;
        RECT 0.060 2090.730 2956.180 2131.630 ;
        RECT 0.060 2045.730 2956.180 2086.630 ;
        RECT 0.060 2000.730 2956.180 2041.630 ;
        RECT 0.060 1955.730 2956.180 1996.630 ;
        RECT 0.060 1910.730 2956.180 1951.630 ;
        RECT 0.060 1865.730 2956.180 1906.630 ;
        RECT 0.060 1820.730 2956.180 1861.630 ;
        RECT 0.060 1775.730 2956.180 1816.630 ;
        RECT 0.060 1730.730 2956.180 1771.630 ;
        RECT 0.060 1685.730 2956.180 1726.630 ;
        RECT 0.060 1640.730 2956.180 1681.630 ;
        RECT 0.060 1595.730 2956.180 1636.630 ;
        RECT 0.060 1550.730 2956.180 1591.630 ;
        RECT 0.060 1505.730 2956.180 1546.630 ;
        RECT 0.060 1460.730 2956.180 1501.630 ;
        RECT 0.060 1415.730 2956.180 1456.630 ;
        RECT 0.060 1370.730 2956.180 1411.630 ;
        RECT 0.060 1325.730 2956.180 1366.630 ;
        RECT 0.060 1280.730 2956.180 1321.630 ;
        RECT 0.060 1235.730 2956.180 1276.630 ;
        RECT 0.060 1190.730 2956.180 1231.630 ;
        RECT 0.060 1145.730 2956.180 1186.630 ;
        RECT 0.060 1100.730 2956.180 1141.630 ;
        RECT 0.060 1055.730 2956.180 1096.630 ;
        RECT 0.060 1010.730 2956.180 1051.630 ;
        RECT 0.060 965.730 2956.180 1006.630 ;
        RECT 0.060 920.730 2956.180 961.630 ;
        RECT 0.060 875.730 2956.180 916.630 ;
        RECT 0.060 830.730 2956.180 871.630 ;
        RECT 0.060 785.730 2956.180 826.630 ;
        RECT 0.060 740.730 2956.180 781.630 ;
        RECT 0.060 695.730 2956.180 736.630 ;
        RECT 0.060 650.730 2956.180 691.630 ;
        RECT 0.060 605.730 2956.180 646.630 ;
        RECT 0.060 560.730 2956.180 601.630 ;
        RECT 736.740 556.630 2901.660 560.730 ;
        RECT 0.060 515.730 2956.180 556.630 ;
        RECT 0.060 470.730 2956.180 511.630 ;
        RECT 0.060 425.730 2956.180 466.630 ;
        RECT 0.060 380.730 2956.180 421.630 ;
        RECT 0.060 335.730 2956.180 376.630 ;
        RECT 0.060 290.730 2956.180 331.630 ;
        RECT 0.060 245.730 2956.180 286.630 ;
        RECT 0.060 200.730 2956.180 241.630 ;
        RECT 0.060 155.730 2956.180 196.630 ;
        RECT 0.060 110.730 2956.180 151.630 ;
        RECT 0.060 65.730 2956.180 106.630 ;
        RECT 0.060 20.730 2956.180 61.630 ;
        RECT 0.060 1.180 2956.180 16.630 ;
  END
END user_project_wrapper
END LIBRARY

