VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_ctrl
  CLASS BLOCK ;
  FOREIGN efuse_ctrl ;
  ORIGIN 0.000 0.000 ;
  SIZE 2175.000 BY 2370.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 25.920 15.380 27.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 15.380 217.520 49.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 788.115 217.520 809.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 1548.115 217.520 1569.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.920 2308.115 217.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 15.380 407.520 52.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 787.505 407.520 812.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 1547.505 407.520 1572.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 405.920 2307.505 407.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 15.380 597.520 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 787.505 597.520 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 1547.505 597.520 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 2307.505 597.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 15.380 787.520 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 787.530 787.520 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 1547.530 787.520 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.920 2307.530 787.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 15.380 977.520 52.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 787.505 977.520 812.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 1547.505 977.520 1572.245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 975.920 2307.505 977.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1165.920 15.380 1167.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1355.920 15.380 1357.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 15.380 1547.520 49.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 787.530 1547.520 809.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 1547.530 1547.520 1569.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.920 2307.530 1547.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 15.380 1737.520 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 787.505 1737.520 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 1547.505 1737.520 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.920 2307.505 1737.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 15.380 1927.520 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 787.505 1927.520 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 1547.505 1927.520 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1925.920 2307.505 1927.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 15.380 2117.520 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 787.530 2117.520 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 1547.530 2117.520 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2115.920 2307.530 2117.520 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 42.820 111.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 803.300 199.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 1563.780 287.800 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 803.300 111.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 42.820 199.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 1563.780 375.720 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 110.360 1563.780 111.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 42.820 287.800 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 803.300 375.720 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.280 1563.780 199.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.200 803.300 287.800 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 42.820 375.720 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.600 42.820 464.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.520 803.300 552.120 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 1563.780 640.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.600 803.300 464.200 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.520 42.820 552.120 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 1563.780 727.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.600 1563.780 464.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 42.820 640.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 803.300 727.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.520 1563.780 552.120 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 638.440 803.300 640.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 726.360 42.820 727.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 42.820 815.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 803.300 903.800 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 995.160 1563.780 996.760 2309.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 803.300 815.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 42.820 903.800 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.600 1563.780 1080.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 1563.780 815.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 995.160 42.820 996.760 788.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.600 803.300 1080.200 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 902.200 1563.780 903.800 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 995.160 803.300 996.760 1548.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1078.600 42.820 1080.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 42.820 1256.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 1563.780 1431.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 803.300 1256.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 1563.780 1519.800 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.440 1563.780 1256.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 42.820 1431.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 803.300 1519.800 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1430.280 803.300 1431.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1518.200 42.820 1519.800 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 42.820 1607.720 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.600 803.300 1696.200 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1782.520 1563.780 1784.120 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 803.300 1607.720 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.600 42.820 1696.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 1563.780 1872.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1606.120 1563.780 1607.720 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1782.520 42.820 1784.120 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 803.300 1872.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1694.600 1563.780 1696.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1782.520 803.300 1784.120 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1870.440 42.820 1872.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 42.820 1959.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 803.300 2047.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2142.600 1563.780 2144.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 803.300 1959.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 42.820 2047.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1958.360 1563.780 1959.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2142.600 42.820 2144.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2046.280 1563.780 2047.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2142.600 803.300 2144.200 1552.620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 35.520 15.380 37.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 15.380 227.120 49.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 787.530 227.120 809.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 1547.530 227.120 1569.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 225.520 2307.530 227.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 15.380 417.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 787.505 417.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 1547.505 417.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.520 2307.505 417.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 15.380 607.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 787.505 607.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 1547.505 607.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.520 2307.505 607.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 15.380 797.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 787.530 797.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 1547.530 797.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 795.520 2307.530 797.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 985.520 15.380 987.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1175.520 15.380 1177.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 15.380 1367.120 49.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 787.530 1367.120 809.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 1547.530 1367.120 1569.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.520 2307.530 1367.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 15.380 1557.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 787.505 1557.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 1547.505 1557.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.520 2307.505 1557.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 15.380 1747.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 787.505 1747.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 1547.505 1747.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1745.520 2307.505 1747.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 15.380 1937.120 52.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 787.530 1937.120 812.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 1547.530 1937.120 1572.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1935.520 2307.530 1937.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 15.380 2127.120 50.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 788.115 2127.120 810.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 1548.115 2127.120 1570.510 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2125.520 2308.115 2127.120 2352.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 42.820 122.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 803.300 209.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 1563.780 297.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 803.300 122.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 42.820 209.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 1563.780 385.800 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.440 1563.780 122.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 42.820 297.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 803.300 385.800 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.360 1563.780 209.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.280 803.300 297.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 384.200 42.820 385.800 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.680 42.820 474.280 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.600 803.300 562.200 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 1563.780 650.120 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.680 803.300 474.280 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.600 42.820 562.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 1563.780 738.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.680 1563.780 474.280 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 42.820 650.120 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 803.300 738.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.600 1563.780 562.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.520 803.300 650.120 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.440 42.820 738.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 42.820 825.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 803.300 913.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 803.300 825.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 42.820 913.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.680 1563.780 1090.280 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 824.360 1563.780 825.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.680 803.300 1090.280 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.280 1563.780 913.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.680 42.820 1090.280 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 42.820 1266.120 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.840 807.220 1348.440 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 1563.780 1441.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 803.300 1266.120 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.840 46.740 1348.440 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 1563.780 1529.880 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.520 1563.780 1266.120 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 42.820 1441.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 803.300 1529.880 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.840 1567.700 1348.440 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.360 803.300 1441.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1528.280 42.820 1529.880 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 42.820 1617.800 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.680 803.300 1706.280 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.600 1563.780 1794.200 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 803.300 1617.800 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.680 42.820 1706.280 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 1563.780 1882.120 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1616.200 1563.780 1617.800 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.600 42.820 1794.200 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 803.300 1882.120 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.680 1563.780 1706.280 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1792.600 803.300 1794.200 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1880.520 42.820 1882.120 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 42.820 1970.040 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 803.300 2057.960 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2152.680 1563.780 2154.280 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 803.300 1970.040 1552.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 42.820 2057.960 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.440 1563.780 1970.040 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2152.680 42.820 2154.280 792.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2056.360 1563.780 2057.960 2313.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2152.680 803.300 2154.280 1552.620 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1884.960 0.000 1885.520 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 0.000 417.200 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 0.000 608.720 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2076.480 0.000 2077.040 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2012.640 0.000 2013.200 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1246.560 0.000 1247.120 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1310.400 0.000 1310.960 4.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 0.000 1374.800 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1438.080 0.000 1438.640 4.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1501.920 0.000 1502.480 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1565.760 0.000 1566.320 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 0.000 1630.160 4.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1693.440 0.000 1694.000 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 0.000 800.240 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 0.000 864.080 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 0.000 927.920 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 0.000 1055.600 4.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 0.000 1119.440 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1182.720 0.000 1183.280 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2140.320 0.000 2140.880 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1948.800 0.000 1949.360 4.000 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1821.120 0.000 1821.680 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 0.000 1757.840 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2167.760 2352.300 ;
      LAYER Metal2 ;
        RECT 24.780 4.300 2154.140 2352.190 ;
        RECT 24.780 3.500 33.300 4.300 ;
        RECT 34.460 3.500 97.140 4.300 ;
        RECT 98.300 3.500 160.980 4.300 ;
        RECT 162.140 3.500 224.820 4.300 ;
        RECT 225.980 3.500 288.660 4.300 ;
        RECT 289.820 3.500 352.500 4.300 ;
        RECT 353.660 3.500 416.340 4.300 ;
        RECT 417.500 3.500 480.180 4.300 ;
        RECT 481.340 3.500 544.020 4.300 ;
        RECT 545.180 3.500 607.860 4.300 ;
        RECT 609.020 3.500 671.700 4.300 ;
        RECT 672.860 3.500 735.540 4.300 ;
        RECT 736.700 3.500 799.380 4.300 ;
        RECT 800.540 3.500 863.220 4.300 ;
        RECT 864.380 3.500 927.060 4.300 ;
        RECT 928.220 3.500 990.900 4.300 ;
        RECT 992.060 3.500 1054.740 4.300 ;
        RECT 1055.900 3.500 1118.580 4.300 ;
        RECT 1119.740 3.500 1182.420 4.300 ;
        RECT 1183.580 3.500 1246.260 4.300 ;
        RECT 1247.420 3.500 1310.100 4.300 ;
        RECT 1311.260 3.500 1373.940 4.300 ;
        RECT 1375.100 3.500 1437.780 4.300 ;
        RECT 1438.940 3.500 1501.620 4.300 ;
        RECT 1502.780 3.500 1565.460 4.300 ;
        RECT 1566.620 3.500 1629.300 4.300 ;
        RECT 1630.460 3.500 1693.140 4.300 ;
        RECT 1694.300 3.500 1756.980 4.300 ;
        RECT 1758.140 3.500 1820.820 4.300 ;
        RECT 1821.980 3.500 1884.660 4.300 ;
        RECT 1885.820 3.500 1948.500 4.300 ;
        RECT 1949.660 3.500 2012.340 4.300 ;
        RECT 2013.500 3.500 2076.180 4.300 ;
        RECT 2077.340 3.500 2140.020 4.300 ;
        RECT 2141.180 3.500 2154.140 4.300 ;
      LAYER Metal3 ;
        RECT 24.170 15.540 2154.190 2352.140 ;
      LAYER Metal4 ;
        RECT 24.220 18.010 25.620 2297.835 ;
        RECT 27.820 18.010 35.220 2297.835 ;
        RECT 37.420 1563.480 110.060 2297.835 ;
        RECT 112.260 1563.480 120.140 2297.835 ;
        RECT 122.340 1563.480 197.980 2297.835 ;
        RECT 200.180 1563.480 208.060 2297.835 ;
        RECT 210.260 1570.020 285.900 2297.835 ;
        RECT 210.260 1563.480 215.620 1570.020 ;
        RECT 37.420 1552.920 215.620 1563.480 ;
        RECT 37.420 803.000 110.060 1552.920 ;
        RECT 112.260 803.000 120.140 1552.920 ;
        RECT 122.340 803.000 197.980 1552.920 ;
        RECT 200.180 803.000 208.060 1552.920 ;
        RECT 210.260 1547.815 215.620 1552.920 ;
        RECT 217.820 1547.815 225.220 1570.020 ;
        RECT 210.260 1547.230 225.220 1547.815 ;
        RECT 227.420 1563.480 285.900 1570.020 ;
        RECT 288.100 1563.480 295.980 2297.835 ;
        RECT 298.180 1563.480 373.820 2297.835 ;
        RECT 376.020 1563.480 383.900 2297.835 ;
        RECT 386.100 1572.570 462.300 2297.835 ;
        RECT 386.100 1572.545 415.220 1572.570 ;
        RECT 386.100 1563.480 405.620 1572.545 ;
        RECT 227.420 1552.920 405.620 1563.480 ;
        RECT 227.420 1547.230 285.900 1552.920 ;
        RECT 210.260 810.020 285.900 1547.230 ;
        RECT 210.260 803.000 215.620 810.020 ;
        RECT 37.420 792.440 215.620 803.000 ;
        RECT 37.420 42.520 110.060 792.440 ;
        RECT 112.260 42.520 120.140 792.440 ;
        RECT 122.340 42.520 197.980 792.440 ;
        RECT 200.180 42.520 208.060 792.440 ;
        RECT 210.260 787.815 215.620 792.440 ;
        RECT 217.820 787.815 225.220 810.020 ;
        RECT 210.260 787.230 225.220 787.815 ;
        RECT 227.420 803.000 285.900 810.020 ;
        RECT 288.100 803.000 295.980 1552.920 ;
        RECT 298.180 803.000 373.820 1552.920 ;
        RECT 376.020 803.000 383.900 1552.920 ;
        RECT 386.100 1547.205 405.620 1552.920 ;
        RECT 407.820 1547.205 415.220 1572.545 ;
        RECT 417.420 1563.480 462.300 1572.570 ;
        RECT 464.500 1563.480 472.380 2297.835 ;
        RECT 474.580 1563.480 550.220 2297.835 ;
        RECT 552.420 1563.480 560.300 2297.835 ;
        RECT 562.500 1572.570 638.140 2297.835 ;
        RECT 562.500 1563.480 595.620 1572.570 ;
        RECT 417.420 1552.920 595.620 1563.480 ;
        RECT 417.420 1547.205 462.300 1552.920 ;
        RECT 386.100 812.570 462.300 1547.205 ;
        RECT 386.100 812.545 415.220 812.570 ;
        RECT 386.100 803.000 405.620 812.545 ;
        RECT 227.420 792.440 405.620 803.000 ;
        RECT 227.420 787.230 285.900 792.440 ;
        RECT 210.260 50.020 285.900 787.230 ;
        RECT 210.260 42.520 215.620 50.020 ;
        RECT 37.420 18.010 215.620 42.520 ;
        RECT 217.820 18.010 225.220 50.020 ;
        RECT 227.420 42.520 285.900 50.020 ;
        RECT 288.100 42.520 295.980 792.440 ;
        RECT 298.180 42.520 373.820 792.440 ;
        RECT 376.020 42.520 383.900 792.440 ;
        RECT 386.100 787.205 405.620 792.440 ;
        RECT 407.820 787.205 415.220 812.545 ;
        RECT 417.420 803.000 462.300 812.570 ;
        RECT 464.500 803.000 472.380 1552.920 ;
        RECT 474.580 803.000 550.220 1552.920 ;
        RECT 552.420 803.000 560.300 1552.920 ;
        RECT 562.500 1547.205 595.620 1552.920 ;
        RECT 597.820 1547.205 605.220 1572.570 ;
        RECT 607.420 1563.480 638.140 1572.570 ;
        RECT 640.340 1563.480 648.220 2297.835 ;
        RECT 650.420 1563.480 726.060 2297.835 ;
        RECT 728.260 1563.480 736.140 2297.835 ;
        RECT 738.340 1572.570 813.980 2297.835 ;
        RECT 738.340 1563.480 785.620 1572.570 ;
        RECT 607.420 1552.920 785.620 1563.480 ;
        RECT 607.420 1547.205 638.140 1552.920 ;
        RECT 562.500 812.570 638.140 1547.205 ;
        RECT 562.500 803.000 595.620 812.570 ;
        RECT 417.420 792.440 595.620 803.000 ;
        RECT 417.420 787.205 462.300 792.440 ;
        RECT 386.100 52.570 462.300 787.205 ;
        RECT 386.100 52.545 415.220 52.570 ;
        RECT 386.100 42.520 405.620 52.545 ;
        RECT 227.420 18.010 405.620 42.520 ;
        RECT 407.820 18.010 415.220 52.545 ;
        RECT 417.420 42.520 462.300 52.570 ;
        RECT 464.500 42.520 472.380 792.440 ;
        RECT 474.580 42.520 550.220 792.440 ;
        RECT 552.420 42.520 560.300 792.440 ;
        RECT 562.500 787.205 595.620 792.440 ;
        RECT 597.820 787.205 605.220 812.570 ;
        RECT 607.420 803.000 638.140 812.570 ;
        RECT 640.340 803.000 648.220 1552.920 ;
        RECT 650.420 803.000 726.060 1552.920 ;
        RECT 728.260 803.000 736.140 1552.920 ;
        RECT 738.340 1547.230 785.620 1552.920 ;
        RECT 787.820 1547.230 795.220 1572.570 ;
        RECT 797.420 1563.480 813.980 1572.570 ;
        RECT 816.180 1563.480 824.060 2297.835 ;
        RECT 826.260 1563.480 901.900 2297.835 ;
        RECT 904.100 1563.480 911.980 2297.835 ;
        RECT 914.180 1572.545 985.220 2297.835 ;
        RECT 914.180 1563.480 975.620 1572.545 ;
        RECT 797.420 1552.920 975.620 1563.480 ;
        RECT 797.420 1547.230 813.980 1552.920 ;
        RECT 738.340 812.570 813.980 1547.230 ;
        RECT 738.340 803.000 785.620 812.570 ;
        RECT 607.420 792.440 785.620 803.000 ;
        RECT 607.420 787.205 638.140 792.440 ;
        RECT 562.500 52.570 638.140 787.205 ;
        RECT 562.500 42.520 595.620 52.570 ;
        RECT 417.420 18.010 595.620 42.520 ;
        RECT 597.820 18.010 605.220 52.570 ;
        RECT 607.420 42.520 638.140 52.570 ;
        RECT 640.340 42.520 648.220 792.440 ;
        RECT 650.420 42.520 726.060 792.440 ;
        RECT 728.260 42.520 736.140 792.440 ;
        RECT 738.340 787.230 785.620 792.440 ;
        RECT 787.820 787.230 795.220 812.570 ;
        RECT 797.420 803.000 813.980 812.570 ;
        RECT 816.180 803.000 824.060 1552.920 ;
        RECT 826.260 803.000 901.900 1552.920 ;
        RECT 904.100 803.000 911.980 1552.920 ;
        RECT 914.180 1547.205 975.620 1552.920 ;
        RECT 977.820 1547.205 985.220 1572.545 ;
        RECT 914.180 812.545 985.220 1547.205 ;
        RECT 914.180 803.000 975.620 812.545 ;
        RECT 797.420 792.440 975.620 803.000 ;
        RECT 797.420 787.230 813.980 792.440 ;
        RECT 738.340 52.570 813.980 787.230 ;
        RECT 738.340 42.520 785.620 52.570 ;
        RECT 607.420 18.010 785.620 42.520 ;
        RECT 787.820 18.010 795.220 52.570 ;
        RECT 797.420 42.520 813.980 52.570 ;
        RECT 816.180 42.520 824.060 792.440 ;
        RECT 826.260 42.520 901.900 792.440 ;
        RECT 904.100 42.520 911.980 792.440 ;
        RECT 914.180 787.205 975.620 792.440 ;
        RECT 977.820 787.205 985.220 812.545 ;
        RECT 914.180 52.545 985.220 787.205 ;
        RECT 914.180 42.520 975.620 52.545 ;
        RECT 797.420 18.010 975.620 42.520 ;
        RECT 977.820 18.010 985.220 52.545 ;
        RECT 987.420 1563.480 994.860 2297.835 ;
        RECT 997.060 1563.480 1078.300 2297.835 ;
        RECT 1080.500 1563.480 1088.380 2297.835 ;
        RECT 1090.580 1563.480 1165.620 2297.835 ;
        RECT 987.420 1552.920 1165.620 1563.480 ;
        RECT 987.420 1549.000 1078.300 1552.920 ;
        RECT 987.420 803.000 994.860 1549.000 ;
        RECT 997.060 803.000 1078.300 1549.000 ;
        RECT 1080.500 803.000 1088.380 1552.920 ;
        RECT 1090.580 803.000 1165.620 1552.920 ;
        RECT 987.420 792.440 1165.620 803.000 ;
        RECT 987.420 788.520 1078.300 792.440 ;
        RECT 987.420 42.520 994.860 788.520 ;
        RECT 997.060 42.520 1078.300 788.520 ;
        RECT 1080.500 42.520 1088.380 792.440 ;
        RECT 1090.580 42.520 1165.620 792.440 ;
        RECT 987.420 18.010 1165.620 42.520 ;
        RECT 1167.820 18.010 1175.220 2297.835 ;
        RECT 1177.420 1563.480 1254.140 2297.835 ;
        RECT 1256.340 1563.480 1264.220 2297.835 ;
        RECT 1266.420 1567.400 1346.540 2297.835 ;
        RECT 1348.740 1567.400 1355.620 2297.835 ;
        RECT 1266.420 1563.480 1355.620 1567.400 ;
        RECT 1177.420 1552.920 1355.620 1563.480 ;
        RECT 1177.420 803.000 1254.140 1552.920 ;
        RECT 1256.340 803.000 1264.220 1552.920 ;
        RECT 1266.420 806.920 1346.540 1552.920 ;
        RECT 1348.740 806.920 1355.620 1552.920 ;
        RECT 1266.420 803.000 1355.620 806.920 ;
        RECT 1177.420 792.440 1355.620 803.000 ;
        RECT 1177.420 42.520 1254.140 792.440 ;
        RECT 1256.340 42.520 1264.220 792.440 ;
        RECT 1266.420 46.440 1346.540 792.440 ;
        RECT 1348.740 46.440 1355.620 792.440 ;
        RECT 1266.420 42.520 1355.620 46.440 ;
        RECT 1177.420 18.010 1355.620 42.520 ;
        RECT 1357.820 1570.020 1429.980 2297.835 ;
        RECT 1357.820 1547.230 1365.220 1570.020 ;
        RECT 1367.420 1563.480 1429.980 1570.020 ;
        RECT 1432.180 1563.480 1440.060 2297.835 ;
        RECT 1442.260 1563.480 1517.900 2297.835 ;
        RECT 1520.100 1563.480 1527.980 2297.835 ;
        RECT 1530.180 1572.570 1605.820 2297.835 ;
        RECT 1530.180 1570.020 1555.220 1572.570 ;
        RECT 1530.180 1563.480 1545.620 1570.020 ;
        RECT 1367.420 1552.920 1545.620 1563.480 ;
        RECT 1367.420 1547.230 1429.980 1552.920 ;
        RECT 1357.820 810.020 1429.980 1547.230 ;
        RECT 1357.820 787.230 1365.220 810.020 ;
        RECT 1367.420 803.000 1429.980 810.020 ;
        RECT 1432.180 803.000 1440.060 1552.920 ;
        RECT 1442.260 803.000 1517.900 1552.920 ;
        RECT 1520.100 803.000 1527.980 1552.920 ;
        RECT 1530.180 1547.230 1545.620 1552.920 ;
        RECT 1547.820 1547.230 1555.220 1570.020 ;
        RECT 1530.180 1547.205 1555.220 1547.230 ;
        RECT 1557.420 1563.480 1605.820 1572.570 ;
        RECT 1608.020 1563.480 1615.900 2297.835 ;
        RECT 1618.100 1563.480 1694.300 2297.835 ;
        RECT 1696.500 1563.480 1704.380 2297.835 ;
        RECT 1706.580 1572.570 1782.220 2297.835 ;
        RECT 1706.580 1563.480 1735.620 1572.570 ;
        RECT 1557.420 1552.920 1735.620 1563.480 ;
        RECT 1557.420 1547.205 1605.820 1552.920 ;
        RECT 1530.180 812.570 1605.820 1547.205 ;
        RECT 1530.180 810.020 1555.220 812.570 ;
        RECT 1530.180 803.000 1545.620 810.020 ;
        RECT 1367.420 792.440 1545.620 803.000 ;
        RECT 1367.420 787.230 1429.980 792.440 ;
        RECT 1357.820 50.020 1429.980 787.230 ;
        RECT 1357.820 18.010 1365.220 50.020 ;
        RECT 1367.420 42.520 1429.980 50.020 ;
        RECT 1432.180 42.520 1440.060 792.440 ;
        RECT 1442.260 42.520 1517.900 792.440 ;
        RECT 1520.100 42.520 1527.980 792.440 ;
        RECT 1530.180 787.230 1545.620 792.440 ;
        RECT 1547.820 787.230 1555.220 810.020 ;
        RECT 1530.180 787.205 1555.220 787.230 ;
        RECT 1557.420 803.000 1605.820 812.570 ;
        RECT 1608.020 803.000 1615.900 1552.920 ;
        RECT 1618.100 803.000 1694.300 1552.920 ;
        RECT 1696.500 803.000 1704.380 1552.920 ;
        RECT 1706.580 1547.205 1735.620 1552.920 ;
        RECT 1737.820 1547.205 1745.220 1572.570 ;
        RECT 1747.420 1563.480 1782.220 1572.570 ;
        RECT 1784.420 1563.480 1792.300 2297.835 ;
        RECT 1794.500 1563.480 1870.140 2297.835 ;
        RECT 1872.340 1563.480 1880.220 2297.835 ;
        RECT 1882.420 1572.570 1958.060 2297.835 ;
        RECT 1882.420 1563.480 1925.620 1572.570 ;
        RECT 1747.420 1552.920 1925.620 1563.480 ;
        RECT 1747.420 1547.205 1782.220 1552.920 ;
        RECT 1706.580 812.570 1782.220 1547.205 ;
        RECT 1706.580 803.000 1735.620 812.570 ;
        RECT 1557.420 792.440 1735.620 803.000 ;
        RECT 1557.420 787.205 1605.820 792.440 ;
        RECT 1530.180 52.570 1605.820 787.205 ;
        RECT 1530.180 50.020 1555.220 52.570 ;
        RECT 1530.180 42.520 1545.620 50.020 ;
        RECT 1367.420 18.010 1545.620 42.520 ;
        RECT 1547.820 18.010 1555.220 50.020 ;
        RECT 1557.420 42.520 1605.820 52.570 ;
        RECT 1608.020 42.520 1615.900 792.440 ;
        RECT 1618.100 42.520 1694.300 792.440 ;
        RECT 1696.500 42.520 1704.380 792.440 ;
        RECT 1706.580 787.205 1735.620 792.440 ;
        RECT 1737.820 787.205 1745.220 812.570 ;
        RECT 1747.420 803.000 1782.220 812.570 ;
        RECT 1784.420 803.000 1792.300 1552.920 ;
        RECT 1794.500 803.000 1870.140 1552.920 ;
        RECT 1872.340 803.000 1880.220 1552.920 ;
        RECT 1882.420 1547.205 1925.620 1552.920 ;
        RECT 1927.820 1547.230 1935.220 1572.570 ;
        RECT 1937.420 1563.480 1958.060 1572.570 ;
        RECT 1960.260 1563.480 1968.140 2297.835 ;
        RECT 1970.340 1563.480 2045.980 2297.835 ;
        RECT 2048.180 1563.480 2056.060 2297.835 ;
        RECT 2058.260 1572.570 2134.020 2297.835 ;
        RECT 2058.260 1563.480 2115.620 1572.570 ;
        RECT 1937.420 1552.920 2115.620 1563.480 ;
        RECT 1937.420 1547.230 1958.060 1552.920 ;
        RECT 1927.820 1547.205 1958.060 1547.230 ;
        RECT 1882.420 812.570 1958.060 1547.205 ;
        RECT 1882.420 803.000 1925.620 812.570 ;
        RECT 1747.420 792.440 1925.620 803.000 ;
        RECT 1747.420 787.205 1782.220 792.440 ;
        RECT 1706.580 52.570 1782.220 787.205 ;
        RECT 1706.580 42.520 1735.620 52.570 ;
        RECT 1557.420 18.010 1735.620 42.520 ;
        RECT 1737.820 18.010 1745.220 52.570 ;
        RECT 1747.420 42.520 1782.220 52.570 ;
        RECT 1784.420 42.520 1792.300 792.440 ;
        RECT 1794.500 42.520 1870.140 792.440 ;
        RECT 1872.340 42.520 1880.220 792.440 ;
        RECT 1882.420 787.205 1925.620 792.440 ;
        RECT 1927.820 787.230 1935.220 812.570 ;
        RECT 1937.420 803.000 1958.060 812.570 ;
        RECT 1960.260 803.000 1968.140 1552.920 ;
        RECT 1970.340 803.000 2045.980 1552.920 ;
        RECT 2048.180 803.000 2056.060 1552.920 ;
        RECT 2058.260 1547.230 2115.620 1552.920 ;
        RECT 2117.820 1570.810 2134.020 1572.570 ;
        RECT 2117.820 1547.815 2125.220 1570.810 ;
        RECT 2127.420 1547.815 2134.020 1570.810 ;
        RECT 2117.820 1547.230 2134.020 1547.815 ;
        RECT 2058.260 812.570 2134.020 1547.230 ;
        RECT 2058.260 803.000 2115.620 812.570 ;
        RECT 1937.420 792.440 2115.620 803.000 ;
        RECT 1937.420 787.230 1958.060 792.440 ;
        RECT 1927.820 787.205 1958.060 787.230 ;
        RECT 1882.420 52.570 1958.060 787.205 ;
        RECT 1882.420 42.520 1925.620 52.570 ;
        RECT 1747.420 18.010 1925.620 42.520 ;
        RECT 1927.820 18.010 1935.220 52.570 ;
        RECT 1937.420 42.520 1958.060 52.570 ;
        RECT 1960.260 42.520 1968.140 792.440 ;
        RECT 1970.340 42.520 2045.980 792.440 ;
        RECT 2048.180 42.520 2056.060 792.440 ;
        RECT 2058.260 787.230 2115.620 792.440 ;
        RECT 2117.820 810.810 2134.020 812.570 ;
        RECT 2117.820 787.815 2125.220 810.810 ;
        RECT 2127.420 787.815 2134.020 810.810 ;
        RECT 2117.820 787.230 2134.020 787.815 ;
        RECT 2058.260 52.570 2134.020 787.230 ;
        RECT 2058.260 42.520 2115.620 52.570 ;
        RECT 1937.420 18.010 2115.620 42.520 ;
        RECT 2117.820 50.810 2134.020 52.570 ;
        RECT 2117.820 18.010 2125.220 50.810 ;
        RECT 2127.420 18.010 2134.020 50.810 ;
      LAYER Metal5 ;
        RECT 10 0 2165 34.5 ;
        RECT 10 49.5 2165 79.5 ;
        RECT 10 94.5 2165 124.5 ;
        RECT 10 139.5 2165 169.5 ;
        RECT 10 184.5 2165 214.5 ;
        RECT 10 229.5 2165 259.5 ;
        RECT 10 274.5 2165 304.5 ;
        RECT 10 319.5 2165 349.5 ;
        RECT 10 364.5 2165 394.5 ;
        RECT 10 409.5 2165 439.5 ;
        RECT 10 454.5 2165 484.5 ;
        RECT 10 499.5 2165 529.5 ;
        RECT 10 544.5 2165 574.5 ;
        RECT 10 589.5 2165 619.5 ;
        RECT 10 634.5 2165 664.5 ;
        RECT 10 679.5 2165 709.5 ;
        RECT 10 724.5 2165 754.5 ;
        RECT 10 769.5 2165 799.5 ;
        RECT 10 814.5 2165 844.5 ;
        RECT 10 859.5 2165 889.5 ;
        RECT 10 904.5 2165 934.5 ;
        RECT 10 949.5 2165 979.5 ;
        RECT 10 994.5 2165 1024.5 ;
        RECT 10 1039.5 2165 1069.5 ;
        RECT 10 1084.5 2165 1114.5 ;
        RECT 10 1129.5 2165 1159.5 ;
        RECT 10 1174.5 2165 1204.5 ;
        RECT 10 1219.5 2165 1249.5 ;
        RECT 10 1264.5 2165 1294.5 ;
        RECT 10 1309.5 2165 1339.5 ;
        RECT 10 1354.5 2165 1384.5 ;
        RECT 10 1399.5 2165 1429.5 ;
        RECT 10 1444.5 2165 1474.5 ;
        RECT 10 1489.5 2165 1519.5 ;
        RECT 10 1534.5 2165 1564.5 ;
        RECT 10 1579.5 2165 1609.5 ;
        RECT 10 1624.5 2165 1654.5 ;
        RECT 10 1669.5 2165 1699.5 ;
        RECT 10 1714.5 2165 1744.5 ;
        RECT 10 1759.5 2165 1789.5 ;
        RECT 10 1804.5 2165 1834.5 ;
        RECT 10 1849.5 2165 1879.5 ;
        RECT 10 1894.5 2165 1924.5 ;
        RECT 10 1939.5 2165 1969.5 ;
        RECT 10 1984.5 2165 2014.5 ;
        RECT 10 2029.5 2165 2059.5 ;
        RECT 10 2074.5 2165 2104.5 ;
        RECT 10 2119.5 2165 2149.5 ;
        RECT 10 2164.5 2165 2194.5 ;
        RECT 10 2209.5 2165 2239.5 ;
        RECT 10 2254.5 2165 2284.5 ;
        RECT 10 2299.5 2165 2329.5 ;
  END
END efuse_ctrl
END LIBRARY

