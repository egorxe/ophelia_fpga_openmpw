VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_struct_block
  CLASS BLOCK ;
  FOREIGN fpga_struct_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 310.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 16.640 7.540 18.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.640 7.540 68.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.640 7.540 118.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.640 7.540 168.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.640 7.540 218.240 302.140 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 41.640 7.540 43.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 91.640 7.540 93.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 141.640 7.540 143.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 191.640 7.540 193.240 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 241.640 7.540 243.240 302.140 ;
    END
  END VSS
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 11.760 250.000 12.320 ;
    END
  END clk_i
  PIN config_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.640 306.000 11.200 310.000 ;
    END
  END config_clk_i
  PIN config_ena_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 306.000 17.360 310.000 ;
    END
  END config_ena_i
  PIN config_shift_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 306.000 23.520 310.000 ;
    END
  END config_shift_i
  PIN config_shift_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END config_shift_o
  PIN glb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 306.000 29.680 310.000 ;
    END
  END glb_rstn_i
  PIN inputs_down_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END inputs_down_i[0]
  PIN inputs_down_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END inputs_down_i[10]
  PIN inputs_down_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END inputs_down_i[11]
  PIN inputs_down_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END inputs_down_i[12]
  PIN inputs_down_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END inputs_down_i[13]
  PIN inputs_down_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END inputs_down_i[14]
  PIN inputs_down_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END inputs_down_i[15]
  PIN inputs_down_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END inputs_down_i[16]
  PIN inputs_down_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END inputs_down_i[17]
  PIN inputs_down_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END inputs_down_i[18]
  PIN inputs_down_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END inputs_down_i[19]
  PIN inputs_down_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END inputs_down_i[1]
  PIN inputs_down_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END inputs_down_i[20]
  PIN inputs_down_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END inputs_down_i[21]
  PIN inputs_down_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END inputs_down_i[22]
  PIN inputs_down_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END inputs_down_i[23]
  PIN inputs_down_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END inputs_down_i[24]
  PIN inputs_down_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END inputs_down_i[25]
  PIN inputs_down_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END inputs_down_i[26]
  PIN inputs_down_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END inputs_down_i[27]
  PIN inputs_down_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END inputs_down_i[28]
  PIN inputs_down_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END inputs_down_i[29]
  PIN inputs_down_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END inputs_down_i[2]
  PIN inputs_down_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END inputs_down_i[30]
  PIN inputs_down_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END inputs_down_i[31]
  PIN inputs_down_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END inputs_down_i[3]
  PIN inputs_down_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END inputs_down_i[4]
  PIN inputs_down_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END inputs_down_i[5]
  PIN inputs_down_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END inputs_down_i[6]
  PIN inputs_down_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END inputs_down_i[7]
  PIN inputs_down_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END inputs_down_i[8]
  PIN inputs_down_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END inputs_down_i[9]
  PIN inputs_left_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END inputs_left_i[0]
  PIN inputs_left_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END inputs_left_i[10]
  PIN inputs_left_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END inputs_left_i[11]
  PIN inputs_left_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END inputs_left_i[12]
  PIN inputs_left_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END inputs_left_i[13]
  PIN inputs_left_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.080 4.000 150.640 ;
    END
  END inputs_left_i[14]
  PIN inputs_left_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END inputs_left_i[15]
  PIN inputs_left_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END inputs_left_i[16]
  PIN inputs_left_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END inputs_left_i[17]
  PIN inputs_left_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END inputs_left_i[18]
  PIN inputs_left_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END inputs_left_i[19]
  PIN inputs_left_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END inputs_left_i[1]
  PIN inputs_left_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.840 4.000 204.400 ;
    END
  END inputs_left_i[20]
  PIN inputs_left_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END inputs_left_i[21]
  PIN inputs_left_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END inputs_left_i[22]
  PIN inputs_left_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.720 4.000 231.280 ;
    END
  END inputs_left_i[23]
  PIN inputs_left_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 4.000 240.240 ;
    END
  END inputs_left_i[24]
  PIN inputs_left_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.640 4.000 249.200 ;
    END
  END inputs_left_i[25]
  PIN inputs_left_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END inputs_left_i[26]
  PIN inputs_left_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END inputs_left_i[27]
  PIN inputs_left_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END inputs_left_i[28]
  PIN inputs_left_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 284.480 4.000 285.040 ;
    END
  END inputs_left_i[29]
  PIN inputs_left_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END inputs_left_i[2]
  PIN inputs_left_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 293.440 4.000 294.000 ;
    END
  END inputs_left_i[30]
  PIN inputs_left_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END inputs_left_i[31]
  PIN inputs_left_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END inputs_left_i[3]
  PIN inputs_left_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END inputs_left_i[4]
  PIN inputs_left_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 4.000 70.000 ;
    END
  END inputs_left_i[5]
  PIN inputs_left_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END inputs_left_i[6]
  PIN inputs_left_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END inputs_left_i[7]
  PIN inputs_left_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END inputs_left_i[8]
  PIN inputs_left_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END inputs_left_i[9]
  PIN inputs_right_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 36.960 250.000 37.520 ;
    END
  END inputs_right_i[0]
  PIN inputs_right_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 120.960 250.000 121.520 ;
    END
  END inputs_right_i[10]
  PIN inputs_right_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 129.360 250.000 129.920 ;
    END
  END inputs_right_i[11]
  PIN inputs_right_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 137.760 250.000 138.320 ;
    END
  END inputs_right_i[12]
  PIN inputs_right_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 146.160 250.000 146.720 ;
    END
  END inputs_right_i[13]
  PIN inputs_right_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 154.560 250.000 155.120 ;
    END
  END inputs_right_i[14]
  PIN inputs_right_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 162.960 250.000 163.520 ;
    END
  END inputs_right_i[15]
  PIN inputs_right_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 171.360 250.000 171.920 ;
    END
  END inputs_right_i[16]
  PIN inputs_right_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 179.760 250.000 180.320 ;
    END
  END inputs_right_i[17]
  PIN inputs_right_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 188.160 250.000 188.720 ;
    END
  END inputs_right_i[18]
  PIN inputs_right_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 196.560 250.000 197.120 ;
    END
  END inputs_right_i[19]
  PIN inputs_right_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 45.360 250.000 45.920 ;
    END
  END inputs_right_i[1]
  PIN inputs_right_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 204.960 250.000 205.520 ;
    END
  END inputs_right_i[20]
  PIN inputs_right_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 213.360 250.000 213.920 ;
    END
  END inputs_right_i[21]
  PIN inputs_right_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 221.760 250.000 222.320 ;
    END
  END inputs_right_i[22]
  PIN inputs_right_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 230.160 250.000 230.720 ;
    END
  END inputs_right_i[23]
  PIN inputs_right_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 238.560 250.000 239.120 ;
    END
  END inputs_right_i[24]
  PIN inputs_right_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 246.960 250.000 247.520 ;
    END
  END inputs_right_i[25]
  PIN inputs_right_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 255.360 250.000 255.920 ;
    END
  END inputs_right_i[26]
  PIN inputs_right_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 263.760 250.000 264.320 ;
    END
  END inputs_right_i[27]
  PIN inputs_right_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 272.160 250.000 272.720 ;
    END
  END inputs_right_i[28]
  PIN inputs_right_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 280.560 250.000 281.120 ;
    END
  END inputs_right_i[29]
  PIN inputs_right_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 53.760 250.000 54.320 ;
    END
  END inputs_right_i[2]
  PIN inputs_right_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 288.960 250.000 289.520 ;
    END
  END inputs_right_i[30]
  PIN inputs_right_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 297.360 250.000 297.920 ;
    END
  END inputs_right_i[31]
  PIN inputs_right_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 62.160 250.000 62.720 ;
    END
  END inputs_right_i[3]
  PIN inputs_right_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 70.560 250.000 71.120 ;
    END
  END inputs_right_i[4]
  PIN inputs_right_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 78.960 250.000 79.520 ;
    END
  END inputs_right_i[5]
  PIN inputs_right_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 87.360 250.000 87.920 ;
    END
  END inputs_right_i[6]
  PIN inputs_right_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 95.760 250.000 96.320 ;
    END
  END inputs_right_i[7]
  PIN inputs_right_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 104.160 250.000 104.720 ;
    END
  END inputs_right_i[8]
  PIN inputs_right_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 112.560 250.000 113.120 ;
    END
  END inputs_right_i[9]
  PIN inputs_up_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.600 306.000 48.160 310.000 ;
    END
  END inputs_up_i[0]
  PIN inputs_up_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.200 306.000 109.760 310.000 ;
    END
  END inputs_up_i[10]
  PIN inputs_up_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 306.000 115.920 310.000 ;
    END
  END inputs_up_i[11]
  PIN inputs_up_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.520 306.000 122.080 310.000 ;
    END
  END inputs_up_i[12]
  PIN inputs_up_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 306.000 128.240 310.000 ;
    END
  END inputs_up_i[13]
  PIN inputs_up_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.840 306.000 134.400 310.000 ;
    END
  END inputs_up_i[14]
  PIN inputs_up_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 306.000 140.560 310.000 ;
    END
  END inputs_up_i[15]
  PIN inputs_up_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.160 306.000 146.720 310.000 ;
    END
  END inputs_up_i[16]
  PIN inputs_up_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 306.000 152.880 310.000 ;
    END
  END inputs_up_i[17]
  PIN inputs_up_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.480 306.000 159.040 310.000 ;
    END
  END inputs_up_i[18]
  PIN inputs_up_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 306.000 165.200 310.000 ;
    END
  END inputs_up_i[19]
  PIN inputs_up_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 306.000 54.320 310.000 ;
    END
  END inputs_up_i[1]
  PIN inputs_up_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 306.000 171.360 310.000 ;
    END
  END inputs_up_i[20]
  PIN inputs_up_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 306.000 177.520 310.000 ;
    END
  END inputs_up_i[21]
  PIN inputs_up_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.120 306.000 183.680 310.000 ;
    END
  END inputs_up_i[22]
  PIN inputs_up_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 306.000 189.840 310.000 ;
    END
  END inputs_up_i[23]
  PIN inputs_up_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 195.440 306.000 196.000 310.000 ;
    END
  END inputs_up_i[24]
  PIN inputs_up_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 306.000 202.160 310.000 ;
    END
  END inputs_up_i[25]
  PIN inputs_up_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.760 306.000 208.320 310.000 ;
    END
  END inputs_up_i[26]
  PIN inputs_up_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 306.000 214.480 310.000 ;
    END
  END inputs_up_i[27]
  PIN inputs_up_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.080 306.000 220.640 310.000 ;
    END
  END inputs_up_i[28]
  PIN inputs_up_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 306.000 226.800 310.000 ;
    END
  END inputs_up_i[29]
  PIN inputs_up_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.920 306.000 60.480 310.000 ;
    END
  END inputs_up_i[2]
  PIN inputs_up_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 306.000 232.960 310.000 ;
    END
  END inputs_up_i[30]
  PIN inputs_up_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 306.000 239.120 310.000 ;
    END
  END inputs_up_i[31]
  PIN inputs_up_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 306.000 66.640 310.000 ;
    END
  END inputs_up_i[3]
  PIN inputs_up_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 306.000 72.800 310.000 ;
    END
  END inputs_up_i[4]
  PIN inputs_up_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 306.000 78.960 310.000 ;
    END
  END inputs_up_i[5]
  PIN inputs_up_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 306.000 85.120 310.000 ;
    END
  END inputs_up_i[6]
  PIN inputs_up_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 306.000 91.280 310.000 ;
    END
  END inputs_up_i[7]
  PIN inputs_up_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.880 306.000 97.440 310.000 ;
    END
  END inputs_up_i[8]
  PIN inputs_up_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 306.000 103.600 310.000 ;
    END
  END inputs_up_i[9]
  PIN outputs_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.280 306.000 35.840 310.000 ;
    END
  END outputs_o[0]
  PIN outputs_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 20.160 250.000 20.720 ;
    END
  END outputs_o[1]
  PIN outputs_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END outputs_o[2]
  PIN outputs_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END outputs_o[3]
  PIN outputs_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 306.000 42.000 310.000 ;
    END
  END outputs_o[4]
  PIN outputs_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 28.560 250.000 29.120 ;
    END
  END outputs_o[5]
  PIN outputs_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END outputs_o[6]
  PIN outputs_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 4.000 16.240 ;
    END
  END outputs_o[7]
  OBS
      LAYER Metal1 ;
        RECT 1.120 7.540 248.640 303.370 ;
      LAYER Metal2 ;
        RECT 0.140 305.700 10.340 306.740 ;
        RECT 11.500 305.700 16.500 306.740 ;
        RECT 17.660 305.700 22.660 306.740 ;
        RECT 23.820 305.700 28.820 306.740 ;
        RECT 29.980 305.700 34.980 306.740 ;
        RECT 36.140 305.700 41.140 306.740 ;
        RECT 42.300 305.700 47.300 306.740 ;
        RECT 48.460 305.700 53.460 306.740 ;
        RECT 54.620 305.700 59.620 306.740 ;
        RECT 60.780 305.700 65.780 306.740 ;
        RECT 66.940 305.700 71.940 306.740 ;
        RECT 73.100 305.700 78.100 306.740 ;
        RECT 79.260 305.700 84.260 306.740 ;
        RECT 85.420 305.700 90.420 306.740 ;
        RECT 91.580 305.700 96.580 306.740 ;
        RECT 97.740 305.700 102.740 306.740 ;
        RECT 103.900 305.700 108.900 306.740 ;
        RECT 110.060 305.700 115.060 306.740 ;
        RECT 116.220 305.700 121.220 306.740 ;
        RECT 122.380 305.700 127.380 306.740 ;
        RECT 128.540 305.700 133.540 306.740 ;
        RECT 134.700 305.700 139.700 306.740 ;
        RECT 140.860 305.700 145.860 306.740 ;
        RECT 147.020 305.700 152.020 306.740 ;
        RECT 153.180 305.700 158.180 306.740 ;
        RECT 159.340 305.700 164.340 306.740 ;
        RECT 165.500 305.700 170.500 306.740 ;
        RECT 171.660 305.700 176.660 306.740 ;
        RECT 177.820 305.700 182.820 306.740 ;
        RECT 183.980 305.700 188.980 306.740 ;
        RECT 190.140 305.700 195.140 306.740 ;
        RECT 196.300 305.700 201.300 306.740 ;
        RECT 202.460 305.700 207.460 306.740 ;
        RECT 208.620 305.700 213.620 306.740 ;
        RECT 214.780 305.700 219.780 306.740 ;
        RECT 220.940 305.700 225.940 306.740 ;
        RECT 227.100 305.700 232.100 306.740 ;
        RECT 233.260 305.700 238.260 306.740 ;
        RECT 239.420 305.700 249.620 306.740 ;
        RECT 0.140 4.300 249.620 305.700 ;
        RECT 0.140 0.090 9.780 4.300 ;
        RECT 10.940 0.090 16.500 4.300 ;
        RECT 17.660 0.090 23.220 4.300 ;
        RECT 24.380 0.090 29.940 4.300 ;
        RECT 31.100 0.090 36.660 4.300 ;
        RECT 37.820 0.090 43.380 4.300 ;
        RECT 44.540 0.090 50.100 4.300 ;
        RECT 51.260 0.090 56.820 4.300 ;
        RECT 57.980 0.090 63.540 4.300 ;
        RECT 64.700 0.090 70.260 4.300 ;
        RECT 71.420 0.090 76.980 4.300 ;
        RECT 78.140 0.090 83.700 4.300 ;
        RECT 84.860 0.090 90.420 4.300 ;
        RECT 91.580 0.090 97.140 4.300 ;
        RECT 98.300 0.090 103.860 4.300 ;
        RECT 105.020 0.090 110.580 4.300 ;
        RECT 111.740 0.090 117.300 4.300 ;
        RECT 118.460 0.090 124.020 4.300 ;
        RECT 125.180 0.090 130.740 4.300 ;
        RECT 131.900 0.090 137.460 4.300 ;
        RECT 138.620 0.090 144.180 4.300 ;
        RECT 145.340 0.090 150.900 4.300 ;
        RECT 152.060 0.090 157.620 4.300 ;
        RECT 158.780 0.090 164.340 4.300 ;
        RECT 165.500 0.090 171.060 4.300 ;
        RECT 172.220 0.090 177.780 4.300 ;
        RECT 178.940 0.090 184.500 4.300 ;
        RECT 185.660 0.090 191.220 4.300 ;
        RECT 192.380 0.090 197.940 4.300 ;
        RECT 199.100 0.090 204.660 4.300 ;
        RECT 205.820 0.090 211.380 4.300 ;
        RECT 212.540 0.090 218.100 4.300 ;
        RECT 219.260 0.090 224.820 4.300 ;
        RECT 225.980 0.090 231.540 4.300 ;
        RECT 232.700 0.090 238.260 4.300 ;
        RECT 239.420 0.090 249.620 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 303.260 249.670 305.620 ;
        RECT 4.300 302.100 249.670 303.260 ;
        RECT 0.090 298.220 249.670 302.100 ;
        RECT 0.090 297.060 245.700 298.220 ;
        RECT 0.090 294.300 249.670 297.060 ;
        RECT 4.300 293.140 249.670 294.300 ;
        RECT 0.090 289.820 249.670 293.140 ;
        RECT 0.090 288.660 245.700 289.820 ;
        RECT 0.090 285.340 249.670 288.660 ;
        RECT 4.300 284.180 249.670 285.340 ;
        RECT 0.090 281.420 249.670 284.180 ;
        RECT 0.090 280.260 245.700 281.420 ;
        RECT 0.090 276.380 249.670 280.260 ;
        RECT 4.300 275.220 249.670 276.380 ;
        RECT 0.090 273.020 249.670 275.220 ;
        RECT 0.090 271.860 245.700 273.020 ;
        RECT 0.090 267.420 249.670 271.860 ;
        RECT 4.300 266.260 249.670 267.420 ;
        RECT 0.090 264.620 249.670 266.260 ;
        RECT 0.090 263.460 245.700 264.620 ;
        RECT 0.090 258.460 249.670 263.460 ;
        RECT 4.300 257.300 249.670 258.460 ;
        RECT 0.090 256.220 249.670 257.300 ;
        RECT 0.090 255.060 245.700 256.220 ;
        RECT 0.090 249.500 249.670 255.060 ;
        RECT 4.300 248.340 249.670 249.500 ;
        RECT 0.090 247.820 249.670 248.340 ;
        RECT 0.090 246.660 245.700 247.820 ;
        RECT 0.090 240.540 249.670 246.660 ;
        RECT 4.300 239.420 249.670 240.540 ;
        RECT 4.300 239.380 245.700 239.420 ;
        RECT 0.090 238.260 245.700 239.380 ;
        RECT 0.090 231.580 249.670 238.260 ;
        RECT 4.300 231.020 249.670 231.580 ;
        RECT 4.300 230.420 245.700 231.020 ;
        RECT 0.090 229.860 245.700 230.420 ;
        RECT 0.090 222.620 249.670 229.860 ;
        RECT 4.300 221.460 245.700 222.620 ;
        RECT 0.090 214.220 249.670 221.460 ;
        RECT 0.090 213.660 245.700 214.220 ;
        RECT 4.300 213.060 245.700 213.660 ;
        RECT 4.300 212.500 249.670 213.060 ;
        RECT 0.090 205.820 249.670 212.500 ;
        RECT 0.090 204.700 245.700 205.820 ;
        RECT 4.300 204.660 245.700 204.700 ;
        RECT 4.300 203.540 249.670 204.660 ;
        RECT 0.090 197.420 249.670 203.540 ;
        RECT 0.090 196.260 245.700 197.420 ;
        RECT 0.090 195.740 249.670 196.260 ;
        RECT 4.300 194.580 249.670 195.740 ;
        RECT 0.090 189.020 249.670 194.580 ;
        RECT 0.090 187.860 245.700 189.020 ;
        RECT 0.090 186.780 249.670 187.860 ;
        RECT 4.300 185.620 249.670 186.780 ;
        RECT 0.090 180.620 249.670 185.620 ;
        RECT 0.090 179.460 245.700 180.620 ;
        RECT 0.090 177.820 249.670 179.460 ;
        RECT 4.300 176.660 249.670 177.820 ;
        RECT 0.090 172.220 249.670 176.660 ;
        RECT 0.090 171.060 245.700 172.220 ;
        RECT 0.090 168.860 249.670 171.060 ;
        RECT 4.300 167.700 249.670 168.860 ;
        RECT 0.090 163.820 249.670 167.700 ;
        RECT 0.090 162.660 245.700 163.820 ;
        RECT 0.090 159.900 249.670 162.660 ;
        RECT 4.300 158.740 249.670 159.900 ;
        RECT 0.090 155.420 249.670 158.740 ;
        RECT 0.090 154.260 245.700 155.420 ;
        RECT 0.090 150.940 249.670 154.260 ;
        RECT 4.300 149.780 249.670 150.940 ;
        RECT 0.090 147.020 249.670 149.780 ;
        RECT 0.090 145.860 245.700 147.020 ;
        RECT 0.090 141.980 249.670 145.860 ;
        RECT 4.300 140.820 249.670 141.980 ;
        RECT 0.090 138.620 249.670 140.820 ;
        RECT 0.090 137.460 245.700 138.620 ;
        RECT 0.090 133.020 249.670 137.460 ;
        RECT 4.300 131.860 249.670 133.020 ;
        RECT 0.090 130.220 249.670 131.860 ;
        RECT 0.090 129.060 245.700 130.220 ;
        RECT 0.090 124.060 249.670 129.060 ;
        RECT 4.300 122.900 249.670 124.060 ;
        RECT 0.090 121.820 249.670 122.900 ;
        RECT 0.090 120.660 245.700 121.820 ;
        RECT 0.090 115.100 249.670 120.660 ;
        RECT 4.300 113.940 249.670 115.100 ;
        RECT 0.090 113.420 249.670 113.940 ;
        RECT 0.090 112.260 245.700 113.420 ;
        RECT 0.090 106.140 249.670 112.260 ;
        RECT 4.300 105.020 249.670 106.140 ;
        RECT 4.300 104.980 245.700 105.020 ;
        RECT 0.090 103.860 245.700 104.980 ;
        RECT 0.090 97.180 249.670 103.860 ;
        RECT 4.300 96.620 249.670 97.180 ;
        RECT 4.300 96.020 245.700 96.620 ;
        RECT 0.090 95.460 245.700 96.020 ;
        RECT 0.090 88.220 249.670 95.460 ;
        RECT 4.300 87.060 245.700 88.220 ;
        RECT 0.090 79.820 249.670 87.060 ;
        RECT 0.090 79.260 245.700 79.820 ;
        RECT 4.300 78.660 245.700 79.260 ;
        RECT 4.300 78.100 249.670 78.660 ;
        RECT 0.090 71.420 249.670 78.100 ;
        RECT 0.090 70.300 245.700 71.420 ;
        RECT 4.300 70.260 245.700 70.300 ;
        RECT 4.300 69.140 249.670 70.260 ;
        RECT 0.090 63.020 249.670 69.140 ;
        RECT 0.090 61.860 245.700 63.020 ;
        RECT 0.090 61.340 249.670 61.860 ;
        RECT 4.300 60.180 249.670 61.340 ;
        RECT 0.090 54.620 249.670 60.180 ;
        RECT 0.090 53.460 245.700 54.620 ;
        RECT 0.090 52.380 249.670 53.460 ;
        RECT 4.300 51.220 249.670 52.380 ;
        RECT 0.090 46.220 249.670 51.220 ;
        RECT 0.090 45.060 245.700 46.220 ;
        RECT 0.090 43.420 249.670 45.060 ;
        RECT 4.300 42.260 249.670 43.420 ;
        RECT 0.090 37.820 249.670 42.260 ;
        RECT 0.090 36.660 245.700 37.820 ;
        RECT 0.090 34.460 249.670 36.660 ;
        RECT 4.300 33.300 249.670 34.460 ;
        RECT 0.090 29.420 249.670 33.300 ;
        RECT 0.090 28.260 245.700 29.420 ;
        RECT 0.090 25.500 249.670 28.260 ;
        RECT 4.300 24.340 249.670 25.500 ;
        RECT 0.090 21.020 249.670 24.340 ;
        RECT 0.090 19.860 245.700 21.020 ;
        RECT 0.090 16.540 249.670 19.860 ;
        RECT 4.300 15.380 249.670 16.540 ;
        RECT 0.090 12.620 249.670 15.380 ;
        RECT 0.090 11.460 245.700 12.620 ;
        RECT 0.090 7.580 249.670 11.460 ;
        RECT 4.300 6.420 249.670 7.580 ;
        RECT 0.090 0.140 249.670 6.420 ;
      LAYER Metal4 ;
        RECT 4.060 302.440 249.620 305.670 ;
        RECT 4.060 7.240 16.340 302.440 ;
        RECT 18.540 7.240 41.340 302.440 ;
        RECT 43.540 7.240 66.340 302.440 ;
        RECT 68.540 7.240 91.340 302.440 ;
        RECT 93.540 7.240 116.340 302.440 ;
        RECT 118.540 7.240 141.340 302.440 ;
        RECT 143.540 7.240 166.340 302.440 ;
        RECT 168.540 7.240 191.340 302.440 ;
        RECT 193.540 7.240 216.340 302.440 ;
        RECT 218.540 7.240 241.340 302.440 ;
        RECT 243.540 7.240 249.620 302.440 ;
        RECT 4.060 6.250 249.620 7.240 ;
  END
END fpga_struct_block
END LIBRARY

